
module SerialFlashLoader (
	noe_in);	

	input		noe_in;
endmodule
