// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "03/31/2019 11:02:17"

// 
// Device: Altera 5CGXFC5C6F27C6 Package FBGA672
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module SerialFlashLoader (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	noe_in)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	noe_in;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \serial_flash_loader_0|altserial_flash_loader_component|ENHANCED_PGM_QUAD:sfl_inst_enhanced|adapted_tdo~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \noe_in~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \~VCC~combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


SerialFlashLoader_altera_serial_flash_loader serial_flash_loader_0(
	.adapted_tdo(\serial_flash_loader_0|altserial_flash_loader_component|ENHANCED_PGM_QUAD:sfl_inst_enhanced|adapted_tdo~15_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][4]~q ),
	.irf_reg_5_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][5]~q ),
	.irf_reg_6_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][6]~q ),
	.irf_reg_7_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][7]~q ),
	.irf_reg_8_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][8]~q ),
	.irf_reg_9_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][9]~q ),
	.irf_reg_10_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][10]~q ),
	.irf_reg_11_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][11]~q ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][10] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'hDFD5FFFFDFD5FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \~VCC (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~VCC~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~VCC .extended_lut = "off";
defparam \~VCC .lut_mask = 64'h0000000000000000;
defparam \~VCC .shared_arith = "off";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \~QIC_CREATED_GND~I (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~QIC_CREATED_GND~I .extended_lut = "off";
defparam \~QIC_CREATED_GND~I .lut_mask = 64'h0000000000000000;
defparam \~QIC_CREATED_GND~I .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFFB7FFFFFF7BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3 .lut_mask = 64'h5FFF3FFF5FFF3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0 .lut_mask = 64'h7FFFFFFFDFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~VCC~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~VCC~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[11]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~GND~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[10]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~GND~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[9]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~GND~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[8]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~VCC~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[7]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~GND~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~GND~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5 .lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~3_combout ),
	.datab(!\~GND~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~GND~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~VCC~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\~VCC~combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hAAAAAAAAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h55AA55AAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'hAA5555AAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'h66999966FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h96696996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'hF6F9F9F6F6F9F9F6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'hF6F9F9F6F6F9F9F6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'hFEFDFDFEFEFDFDFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'h5F3FFFFF5F3FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\serial_flash_loader_0|altserial_flash_loader_component|ENHANCED_PGM_QUAD:sfl_inst_enhanced|adapted_tdo~15_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'hFAFFFFFFFAFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hEDDEDEEDDEEDEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hFFFFFFFFFDFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hDEDEDEDEDEDEDEDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hDFFFFDFFDFFFFDFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hFFFFD8FFFFFFD8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'hFFF6FFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'hF9F6FFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hFF7FBF3FFF7FBF3F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

assign \noe_in~input_o  = noe_in;

endmodule

module SerialFlashLoader_altera_serial_flash_loader (
	adapted_tdo,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_2,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	irf_reg_5_1,
	irf_reg_6_1,
	irf_reg_7_1,
	irf_reg_8_1,
	irf_reg_9_1,
	irf_reg_10_1,
	irf_reg_11_1)/* synthesis synthesis_greybox=1 */;
output 	adapted_tdo;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_2;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	irf_reg_5_1;
input 	irf_reg_6_1;
input 	irf_reg_7_1;
input 	irf_reg_8_1;
input 	irf_reg_9_1;
input 	irf_reg_10_1;
input 	irf_reg_11_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



SerialFlashLoader_altserial_flash_loader altserial_flash_loader_component(
	.adapted_tdo(adapted_tdo),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_2(state_2),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.irf_reg_5_1(irf_reg_5_1),
	.irf_reg_6_1(irf_reg_6_1),
	.irf_reg_7_1(irf_reg_7_1),
	.irf_reg_8_1(irf_reg_8_1),
	.irf_reg_9_1(irf_reg_9_1),
	.irf_reg_10_1(irf_reg_10_1),
	.irf_reg_11_1(irf_reg_11_1));

endmodule

module SerialFlashLoader_altserial_flash_loader (
	adapted_tdo,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_2,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	irf_reg_5_1,
	irf_reg_6_1,
	irf_reg_7_1,
	irf_reg_8_1,
	irf_reg_9_1,
	irf_reg_10_1,
	irf_reg_11_1)/* synthesis synthesis_greybox=1 */;
output 	adapted_tdo;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_2;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	irf_reg_5_1;
input 	irf_reg_6_1;
input 	irf_reg_7_1;
input 	irf_reg_8_1;
input 	irf_reg_9_1;
input 	irf_reg_10_1;
input 	irf_reg_11_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire data1out_int;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|Equal26~1_combout ;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|single_scein~q ;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|sdoin~reg0_q ;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|data1in~0_combout ;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|data2in~0_combout ;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|data3in~0_combout ;
wire \ENHANCED_PGM_QUAD:sfl_inst_enhanced|dclkin~0_combout ;


SerialFlashLoader_alt_sfl_enhanced_1 \ENHANCED_PGM_QUAD:sfl_inst_enhanced (
	.data1out_int(data1out_int),
	.Equal26(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|Equal26~1_combout ),
	.adapted_tdo(adapted_tdo),
	.single_scein1(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|single_scein~q ),
	.sdoin(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|sdoin~reg0_q ),
	.data1in(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|data1in~0_combout ),
	.data2in(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|data2in~0_combout ),
	.data3in(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|data3in~0_combout ),
	.dclkin(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|dclkin~0_combout ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_2(state_2),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.irf_reg_5_1(irf_reg_5_1),
	.irf_reg_6_1(irf_reg_6_1),
	.irf_reg_7_1(irf_reg_7_1),
	.irf_reg_8_1(irf_reg_8_1),
	.irf_reg_9_1(irf_reg_9_1),
	.irf_reg_10_1(irf_reg_10_1),
	.irf_reg_11_1(irf_reg_11_1));

cyclonev_asmiblock \GEN_ASMI_TYPE_7:asmi_inst (
	.dclk(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|dclkin~0_combout ),
	.sce(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|single_scein~q ),
	.oe(gnd),
	.data0out(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|sdoin~reg0_q ),
	.data1out(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|data1in~0_combout ),
	.data2out(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|data2in~0_combout ),
	.data3out(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|data3in~0_combout ),
	.data0oe(vcc),
	.data1oe(\ENHANCED_PGM_QUAD:sfl_inst_enhanced|Equal26~1_combout ),
	.data2oe(vcc),
	.data3oe(vcc),
	.spidatain(4'b0000),
	.data0in(),
	.data1in(data1out_int),
	.data2in(),
	.data3in(),
	.spisce(),
	.spidclk(),
	.spidataout());
defparam \GEN_ASMI_TYPE_7:asmi_inst .enable_sim = "false";

endmodule

module SerialFlashLoader_alt_sfl_enhanced_1 (
	data1out_int,
	Equal26,
	adapted_tdo,
	single_scein1,
	sdoin,
	data1in,
	data2in,
	data3in,
	dclkin,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_2,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	irf_reg_5_1,
	irf_reg_6_1,
	irf_reg_7_1,
	irf_reg_8_1,
	irf_reg_9_1,
	irf_reg_10_1,
	irf_reg_11_1)/* synthesis synthesis_greybox=1 */;
input 	data1out_int;
output 	Equal26;
output 	adapted_tdo;
output 	single_scein1;
output 	sdoin;
output 	data1in;
output 	data2in;
output 	data3in;
output 	dclkin;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_2;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	irf_reg_5_1;
input 	irf_reg_6_1;
input 	irf_reg_7_1;
input 	irf_reg_8_1;
input 	irf_reg_9_1;
input 	irf_reg_10_1;
input 	irf_reg_11_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_speed_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ;
wire \data_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ;
wire \crc_reg[0]~q ;
wire \crc_reg[1]~q ;
wire \crc_reg[14]~q ;
wire \crc_reg[2]~q ;
wire \crc_reg[13]~q ;
wire \crc_reg[3]~q ;
wire \crc_reg[12]~q ;
wire \crc_reg[4]~q ;
wire \crc_reg[11]~q ;
wire \crc_reg[5]~q ;
wire \crc_reg[10]~q ;
wire \crc_reg[6]~q ;
wire \crc_reg[9]~q ;
wire \crc_reg[7]~q ;
wire \crc_reg[8]~q ;
wire \en4b_reg|dffs[0]~q ;
wire \powerful_reg|dffs[0]~q ;
wire \crc_shifter|dffs[0]~q ;
wire \opcode_reg|dffs[0]~q ;
wire \rstatus_reg|dffs[0]~q ;
wire \rsiid_reg|dffs[0]~q ;
wire \rdi_reg|dffs[0]~q ;
wire \comb~0_combout ;
wire \powerful_reg|dffs[1]~q ;
wire \comb~1_combout ;
wire \reset~q ;
wire \bit_counter|auto_generated|counter_reg_bit[5]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[11]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[10]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[9]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[8]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[7]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[6]~q ;
wire \device_dclk_en_without_sdr~0_combout ;
wire \comb~2_combout ;
wire \bit_counter|auto_generated|counter_reg_bit[4]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[3]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[2]~q ;
wire \bit_counter|auto_generated|counter_reg_bit[1]~q ;
wire \enable_crc_storage~0_combout ;
wire \always5~0_combout ;
wire \comb~3_combout ;
wire \comb~4_combout ;
wire \opcode_reg|dffs[1]~q ;
wire \comb~5_combout ;
wire \comb~6_combout ;
wire \comb~7_combout ;
wire \comb~8_combout ;
wire \comb~9_combout ;
wire \powerful_reg|dffs[2]~q ;
wire \opcode_reg|dffs[7]~q ;
wire \opcode_reg|dffs[6]~q ;
wire \opcode_reg|dffs[5]~q ;
wire \opcode_reg|dffs[4]~q ;
wire \opcode_reg|dffs[2]~q ;
wire \opcode_reg|dffs[3]~q ;
wire \reset_wire~0_combout ;
wire \reset_wire~1_combout ;
wire \sdrs_reg~q ;
wire \comb~11_combout ;
wire \comb~12_combout ;
wire \comb~13_combout ;
wire \powerful_reg|dffs[3]~q ;
wire \crc_shifter_input~0_combout ;
wire \sdrs~combout ;
wire \aai_write_reg|dffs[0]~q ;
wire \aai_data_reg|dffs[0]~q ;
wire \ncso_reg|dffs[0]~q ;
wire \powerful_reg|dffs[4]~q ;
wire \crc_reg[15]~q ;
wire \crc_wire[0]~combout ;
wire \clear_crc~0_combout ;
wire \bit_counter|auto_generated|counter_reg_bit[0]~q ;
wire \clear_crc~1_combout ;
wire \always5~1_combout ;
wire \enable_crc_calculation~0_combout ;
wire \always5~2_combout ;
wire \enable_crc_storage~2_combout ;
wire \enable_crc_change~0_combout ;
wire \crc_reg[14]~0_combout ;
wire \comb~14_combout ;
wire \comb~15_combout ;
wire \comb~16_combout ;
wire \crc_reg~1_combout ;
wire \crc_wire[12]~combout ;
wire \crc_wire[5]~combout ;
wire \Equal11~1_combout ;
wire \Equal5~2_combout ;
wire \Equal26~0_combout ;
wire \Equal17~0_combout ;
wire \Equal11~0_combout ;
wire \Equal6~0_combout ;
wire \Equal14~0_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal10~0_combout ;
wire \Equal6~1_combout ;
wire \Equal3~0_combout ;
wire \Equal16~0_combout ;
wire \Equal16~1_combout ;
wire \Equal15~0_combout ;
wire \Equal11~2_combout ;
wire \adapted_tdo~0_combout ;
wire \Equal3~1_combout ;
wire \Equal3~2_combout ;
wire \Equal5~0_combout ;
wire \adapted_tdo~1_combout ;
wire \adapted_tdo~2_combout ;
wire \Equal5~1_combout ;
wire \Equal5~3_combout ;
wire \bypass_out~q ;
wire \Equal6~2_combout ;
wire \Equal6~3_combout ;
wire \adapted_tdo~3_combout ;
wire \adapted_tdo~4_combout ;
wire \adapted_tdo~5_combout ;
wire \adapted_tdo~6_combout ;
wire \adapted_tdo~7_combout ;
wire \adapted_tdo~8_combout ;
wire \adapted_tdo~9_combout ;
wire \adapted_tdo~10_combout ;
wire \Equal21~0_combout ;
wire \Equal17~1_combout ;
wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \Equal19~0_combout ;
wire \Equal6~4_combout ;
wire \Equal23~0_combout ;
wire \Equal25~0_combout ;
wire \Equal20~0_combout ;
wire \Equal20~1_combout ;
wire \always8~0_combout ;
wire \Equal13~0_combout ;
wire \adapted_tdo~11_combout ;
wire \adapted_tdo~12_combout ;
wire \adapted_tdo~13_combout ;
wire \push_rsiid_inst~0_combout ;
wire \push_rdi_inst~0_combout ;
wire \sdr~combout ;
wire \Equal2~0_combout ;
wire \enable_crc_storage~1_combout ;
wire \LessThan19~0_combout ;
wire \device_dclk_en_without_sdr~1_combout ;
wire \device_dclk_en_without_sdr~2_combout ;
wire \device_dclk_en_without_sdr~3_combout ;
wire \enable_speed_write_data~0_combout ;
wire \always4~0_combout ;
wire \device_dclk_en_without_sdr~4_combout ;
wire \device_dclk_en_without_sdr~5_combout ;
wire \push_rsiid_inst~1_combout ;
wire \always4~1_combout ;
wire \always4~2_combout ;
wire \always4~3_combout ;
wire \LessThan20~0_combout ;
wire \always4~4_combout ;
wire \always4~5_combout ;
wire \device_dclk_en_without_sdr~6_combout ;
wire \Equal23~1_combout ;
wire \always4~6_combout ;
wire \device_dclk_en_without_sdr~7_combout ;
wire \data1out_reg~0_combout ;
wire \data1out_reg~q ;
wire \adapted_tdo~14_combout ;
wire \device_dclk_en_without_sdr~8_combout ;
wire \device_dclk_en_without_sdr~9_combout ;
wire \always4~7_combout ;
wire \always4~8_combout ;
wire \device_dclk_en_without_sdr~10_combout ;
wire \sdoin_wire~0_combout ;
wire \sdoin_wire~1_combout ;
wire \powerful_io0_reg~0_combout ;
wire \udr~combout ;
wire \powerful_ncs_reg~0_combout ;
wire \powerful_io0_reg~q ;
wire \sdoin_wire~3_combout ;
wire \comb~10_combout ;
wire \Equal27~0_combout ;
wire \sdoin_wire~2_combout ;
wire \sdoin_wire~6_combout ;
wire \sdoin_wire~10_combout ;
wire \sdoin_wire~5_combout ;
wire \sdoin_wire~4_combout ;
wire \powerful_io1_reg~0_combout ;
wire \powerful_io1_reg~q ;
wire \powerful_io2_reg~0_combout ;
wire \powerful_io2_reg~q ;
wire \powerful_io3_reg~0_combout ;
wire \powerful_io3_reg~q ;
wire \device_dclk_en_without_sdr~11_combout ;
wire \device_dclk_en~combout ;
wire \device_dclk_en_reg~q ;
wire \powerful_ncs_reg~1_combout ;
wire \powerful_ncs_reg~q ;
wire \udr_reg~q ;
wire \powerful_sck~combout ;
wire \dclkin_without_sdr~combout ;


SerialFlashLoader_lpm_shiftreg_2 aai_write_reg(
	.reset(\reset~q ),
	.dffs_0(\aai_write_reg|dffs[0]~q ),
	.enable(\comb~14_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_10 rdi_reg(
	.dffs_0(\rdi_reg|dffs[0]~q ),
	.reset(\reset~q ),
	.enable(\comb~8_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_11 rsiid_reg(
	.dffs_0(\rsiid_reg|dffs[0]~q ),
	.reset(\reset~q ),
	.enable(\comb~7_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_12 rstatus_reg(
	.dffs_0(\rstatus_reg|dffs[0]~q ),
	.reset(\reset~q ),
	.enable(\comb~6_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_8 opcode_reg(
	.dffs_0(\opcode_reg|dffs[0]~q ),
	.dffs_1(\opcode_reg|dffs[1]~q ),
	.enable(\comb~5_combout ),
	.dffs_7(\opcode_reg|dffs[7]~q ),
	.dffs_6(\opcode_reg|dffs[6]~q ),
	.dffs_5(\opcode_reg|dffs[5]~q ),
	.dffs_4(\opcode_reg|dffs[4]~q ),
	.dffs_2(\opcode_reg|dffs[2]~q ),
	.dffs_3(\opcode_reg|dffs[3]~q ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_counter_1 bit_counter(
	.counter_reg_bit_5(\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.counter_reg_bit_11(\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.counter_reg_bit_10(\bit_counter|auto_generated|counter_reg_bit[10]~q ),
	.counter_reg_bit_9(\bit_counter|auto_generated|counter_reg_bit[9]~q ),
	.counter_reg_bit_8(\bit_counter|auto_generated|counter_reg_bit[8]~q ),
	.counter_reg_bit_7(\bit_counter|auto_generated|counter_reg_bit[7]~q ),
	.counter_reg_bit_6(\bit_counter|auto_generated|counter_reg_bit[6]~q ),
	.counter_reg_bit_4(\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\bit_counter|auto_generated|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\bit_counter|auto_generated|counter_reg_bit[1]~q ),
	.sdrs_reg(\sdrs_reg~q ),
	.comb(\comb~13_combout ),
	.counter_reg_bit_0(\bit_counter|auto_generated|counter_reg_bit[0]~q ),
	.clock(altera_internal_jtag));

SerialFlashLoader_lpm_shiftreg_7 ncso_reg(
	.dffs_0(\ncso_reg|dffs[0]~q ),
	.enable(\comb~16_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_9 powerful_reg(
	.dffs_0(\powerful_reg|dffs[0]~q ),
	.dffs_1(\powerful_reg|dffs[1]~q ),
	.enable(\comb~1_combout ),
	.dffs_2(\powerful_reg|dffs[2]~q ),
	.dffs_3(\powerful_reg|dffs[3]~q ),
	.dffs_4(\powerful_reg|dffs[4]~q ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_3 crc_shifter(
	.dffs_0(\crc_shifter|dffs[0]~q ),
	.reset(\reset~q ),
	.counter_reg_bit_5(\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.device_dclk_en_without_sdr(\device_dclk_en_without_sdr~0_combout ),
	.comb(\comb~2_combout ),
	.enable_crc_storage(\enable_crc_storage~0_combout ),
	.always5(\always5~0_combout ),
	.enable(\comb~3_combout ),
	.crc_shifter_input(\crc_shifter_input~0_combout ),
	.clock(altera_internal_jtag));

SerialFlashLoader_lpm_shiftreg_6 en4b_reg(
	.dffs_0(\en4b_reg|dffs[0]~q ),
	.enable(\comb~0_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_5 data_speed_reg(
	.ram_block8a0(\data_speed_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.Equal3(\Equal3~2_combout ),
	.adapted_tdo(\adapted_tdo~1_combout ),
	.Equal4(\Equal4~1_combout ),
	.sdr(\sdr~combout ),
	.reset(\reset~q ),
	.enable(\comb~4_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_4 data_reg(
	.ram_block8a0(\data_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.Equal19(\Equal19~0_combout ),
	.Equal13(\Equal13~0_combout ),
	.adapted_tdo(\adapted_tdo~11_combout ),
	.sdr(\sdr~combout ),
	.reset(\reset~q ),
	.enable(\comb~9_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

SerialFlashLoader_lpm_shiftreg_1 aai_data_reg(
	.reset(\reset~q ),
	.dffs_0(\aai_data_reg|dffs[0]~q ),
	.enable(\comb~15_combout ),
	.clock(altera_internal_jtag),
	.altera_internal_jtag(altera_internal_jtag1));

dffeas \crc_reg[0] (
	.clk(!altera_internal_jtag),
	.d(\crc_wire[0]~combout ),
	.asdata(\crc_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[0]~q ),
	.prn(vcc));
defparam \crc_reg[0] .is_wysiwyg = "true";
defparam \crc_reg[0] .power_up = "low";

dffeas \crc_reg[1] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[0]~q ),
	.asdata(\crc_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[1]~q ),
	.prn(vcc));
defparam \crc_reg[1] .is_wysiwyg = "true";
defparam \crc_reg[1] .power_up = "low";

dffeas \crc_reg[14] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[13]~q ),
	.asdata(\crc_reg[15]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[14]~q ),
	.prn(vcc));
defparam \crc_reg[14] .is_wysiwyg = "true";
defparam \crc_reg[14] .power_up = "low";

dffeas \crc_reg[2] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[1]~q ),
	.asdata(\crc_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[2]~q ),
	.prn(vcc));
defparam \crc_reg[2] .is_wysiwyg = "true";
defparam \crc_reg[2] .power_up = "low";

dffeas \crc_reg[13] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[12]~q ),
	.asdata(\crc_reg[14]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[13]~q ),
	.prn(vcc));
defparam \crc_reg[13] .is_wysiwyg = "true";
defparam \crc_reg[13] .power_up = "low";

dffeas \crc_reg[3] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[2]~q ),
	.asdata(\crc_reg[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[3]~q ),
	.prn(vcc));
defparam \crc_reg[3] .is_wysiwyg = "true";
defparam \crc_reg[3] .power_up = "low";

dffeas \crc_reg[12] (
	.clk(!altera_internal_jtag),
	.d(\crc_wire[12]~combout ),
	.asdata(\crc_reg[13]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[12]~q ),
	.prn(vcc));
defparam \crc_reg[12] .is_wysiwyg = "true";
defparam \crc_reg[12] .power_up = "low";

dffeas \crc_reg[4] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[3]~q ),
	.asdata(\crc_reg[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[4]~q ),
	.prn(vcc));
defparam \crc_reg[4] .is_wysiwyg = "true";
defparam \crc_reg[4] .power_up = "low";

dffeas \crc_reg[11] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[10]~q ),
	.asdata(\crc_reg[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[11]~q ),
	.prn(vcc));
defparam \crc_reg[11] .is_wysiwyg = "true";
defparam \crc_reg[11] .power_up = "low";

dffeas \crc_reg[5] (
	.clk(!altera_internal_jtag),
	.d(\crc_wire[5]~combout ),
	.asdata(\crc_reg[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[5]~q ),
	.prn(vcc));
defparam \crc_reg[5] .is_wysiwyg = "true";
defparam \crc_reg[5] .power_up = "low";

dffeas \crc_reg[10] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[9]~q ),
	.asdata(\crc_reg[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[10]~q ),
	.prn(vcc));
defparam \crc_reg[10] .is_wysiwyg = "true";
defparam \crc_reg[10] .power_up = "low";

dffeas \crc_reg[6] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[5]~q ),
	.asdata(\crc_reg[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[6]~q ),
	.prn(vcc));
defparam \crc_reg[6] .is_wysiwyg = "true";
defparam \crc_reg[6] .power_up = "low";

dffeas \crc_reg[9] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[8]~q ),
	.asdata(\crc_reg[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[9]~q ),
	.prn(vcc));
defparam \crc_reg[9] .is_wysiwyg = "true";
defparam \crc_reg[9] .power_up = "low";

dffeas \crc_reg[7] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[6]~q ),
	.asdata(\crc_reg[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[7]~q ),
	.prn(vcc));
defparam \crc_reg[7] .is_wysiwyg = "true";
defparam \crc_reg[7] .power_up = "low";

dffeas \crc_reg[8] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg[7]~q ),
	.asdata(\crc_reg[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\always5~1_combout ),
	.sload(\always5~2_combout ),
	.ena(\crc_reg[14]~0_combout ),
	.q(\crc_reg[8]~q ),
	.prn(vcc));
defparam \crc_reg[8] .is_wysiwyg = "true";
defparam \crc_reg[8] .power_up = "low";

cyclonev_lcell_comb \comb~0 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~0_combout ),
	.datac(!\sdr~combout ),
	.datad(!\Equal6~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~1 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\sdr~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~1 .extended_lut = "off";
defparam \comb~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \comb~1 .shared_arith = "off";

dffeas reset(
	.clk(altera_internal_jtag),
	.d(\reset_wire~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset~q ),
	.prn(vcc));
defparam reset.is_wysiwyg = "true";
defparam reset.power_up = "low";

cyclonev_lcell_comb \device_dclk_en_without_sdr~0 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[10]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[9]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[8]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[7]~q ),
	.dataf(!\bit_counter|auto_generated|counter_reg_bit[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~0 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \device_dclk_en_without_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~2 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_5_1),
	.datac(!\Equal5~1_combout ),
	.datad(!\Equal5~2_combout ),
	.datae(!\sdr~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~2 .extended_lut = "off";
defparam \comb~2 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \comb~2 .shared_arith = "off";

cyclonev_lcell_comb \enable_crc_storage~0 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[2]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_crc_storage~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_crc_storage~0 .extended_lut = "off";
defparam \enable_crc_storage~0 .lut_mask = 64'h9669699696696996;
defparam \enable_crc_storage~0 .shared_arith = "off";

cyclonev_lcell_comb \always5~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\Equal1~0_combout ),
	.datac(!\Equal1~1_combout ),
	.datad(!\Equal4~0_combout ),
	.datae(!\sdr~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \always5~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~3 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\device_dclk_en_without_sdr~0_combout ),
	.datac(!\comb~2_combout ),
	.datad(!\enable_crc_storage~0_combout ),
	.datae(!\always5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~3 .extended_lut = "off";
defparam \comb~3 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \comb~3 .shared_arith = "off";

cyclonev_lcell_comb \comb~4 (
	.dataa(!\Equal4~1_combout ),
	.datab(!\Equal3~2_combout ),
	.datac(!\sdr~combout ),
	.datad(!\adapted_tdo~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~4 .extended_lut = "off";
defparam \comb~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \comb~4 .shared_arith = "off";

cyclonev_lcell_comb \comb~5 (
	.dataa(!\Equal10~0_combout ),
	.datab(!\Equal16~1_combout ),
	.datac(!\sdr~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~5 .extended_lut = "off";
defparam \comb~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \comb~5 .shared_arith = "off";

cyclonev_lcell_comb \comb~6 (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal17~0_combout ),
	.datac(!\Equal20~0_combout ),
	.datad(!\Equal11~0_combout ),
	.datae(!\Equal6~0_combout ),
	.dataf(!\sdr~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~6 .extended_lut = "off";
defparam \comb~6 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \comb~6 .shared_arith = "off";

cyclonev_lcell_comb \comb~7 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\Equal21~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(!\Equal15~0_combout ),
	.datae(!\Equal11~2_combout ),
	.dataf(!\sdr~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~7 .extended_lut = "off";
defparam \comb~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \comb~7 .shared_arith = "off";

cyclonev_lcell_comb \comb~8 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\Equal21~0_combout ),
	.datac(!\Equal15~0_combout ),
	.datad(!\sdr~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~8 .extended_lut = "off";
defparam \comb~8 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \comb~8 .shared_arith = "off";

cyclonev_lcell_comb \comb~9 (
	.dataa(!\Equal19~0_combout ),
	.datab(!\Equal13~0_combout ),
	.datac(!\sdr~combout ),
	.datad(!\adapted_tdo~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~9 .extended_lut = "off";
defparam \comb~9 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \comb~9 .shared_arith = "off";

cyclonev_lcell_comb \reset_wire~0 (
	.dataa(!\opcode_reg|dffs[0]~q ),
	.datab(!\opcode_reg|dffs[1]~q ),
	.datac(!\opcode_reg|dffs[2]~q ),
	.datad(!\opcode_reg|dffs[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reset_wire~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reset_wire~0 .extended_lut = "off";
defparam \reset_wire~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \reset_wire~0 .shared_arith = "off";

cyclonev_lcell_comb \reset_wire~1 (
	.dataa(!\sdr~combout ),
	.datab(!\opcode_reg|dffs[7]~q ),
	.datac(!\opcode_reg|dffs[6]~q ),
	.datad(!\opcode_reg|dffs[5]~q ),
	.datae(!\opcode_reg|dffs[4]~q ),
	.dataf(!\reset_wire~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reset_wire~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reset_wire~1 .extended_lut = "off";
defparam \reset_wire~1 .lut_mask = 64'hFFFFFBFFFFFFFFFF;
defparam \reset_wire~1 .shared_arith = "off";

dffeas sdrs_reg(
	.clk(altera_internal_jtag),
	.d(\sdrs~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sdrs_reg~q ),
	.prn(vcc));
defparam sdrs_reg.is_wysiwyg = "true";
defparam sdrs_reg.power_up = "low";

cyclonev_lcell_comb \comb~11 (
	.dataa(!\Equal4~1_combout ),
	.datab(!\Equal20~1_combout ),
	.datac(!\Equal2~0_combout ),
	.datad(!\Equal23~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~11 .extended_lut = "off";
defparam \comb~11 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \comb~11 .shared_arith = "off";

cyclonev_lcell_comb \comb~12 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!state_4),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~12 .extended_lut = "off";
defparam \comb~12 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \comb~12 .shared_arith = "off";

cyclonev_lcell_comb \comb~13 (
	.dataa(!\Equal25~0_combout ),
	.datab(!\Equal5~3_combout ),
	.datac(!\comb~10_combout ),
	.datad(!\comb~11_combout ),
	.datae(!\comb~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~13 .extended_lut = "off";
defparam \comb~13 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \comb~13 .shared_arith = "off";

cyclonev_lcell_comb \crc_shifter_input~0 (
	.dataa(!altera_internal_jtag1),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\device_dclk_en_without_sdr~0_combout ),
	.datad(!\enable_crc_storage~0_combout ),
	.datae(!\always5~0_combout ),
	.dataf(!\crc_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_shifter_input~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_shifter_input~0 .extended_lut = "off";
defparam \crc_shifter_input~0 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \crc_shifter_input~0 .shared_arith = "off";

cyclonev_lcell_comb sdrs(
	.dataa(!virtual_ir_scan_reg),
	.datab(!state_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdrs~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam sdrs.extended_lut = "off";
defparam sdrs.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam sdrs.shared_arith = "off";

dffeas \crc_reg[15] (
	.clk(!altera_internal_jtag),
	.d(\crc_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\crc_reg[15]~q ),
	.prn(vcc));
defparam \crc_reg[15] .is_wysiwyg = "true";
defparam \crc_reg[15] .power_up = "low";

cyclonev_lcell_comb \crc_wire[0] (
	.dataa(!data1out_int),
	.datab(!\crc_reg[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_wire[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_wire[0] .extended_lut = "off";
defparam \crc_wire[0] .lut_mask = 64'h6666666666666666;
defparam \crc_wire[0] .shared_arith = "off";

cyclonev_lcell_comb \clear_crc~0 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clear_crc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \clear_crc~0 .extended_lut = "off";
defparam \clear_crc~0 .lut_mask = 64'h7777777777777777;
defparam \clear_crc~0 .shared_arith = "off";

cyclonev_lcell_comb \clear_crc~1 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[2]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[1]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clear_crc~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \clear_crc~1 .extended_lut = "off";
defparam \clear_crc~1 .lut_mask = 64'hFFFFFF6FFFFFFF6F;
defparam \clear_crc~1 .shared_arith = "off";

cyclonev_lcell_comb \always5~1 (
	.dataa(!\Equal3~2_combout ),
	.datab(!\clear_crc~0_combout ),
	.datac(!\device_dclk_en_without_sdr~0_combout ),
	.datad(!\reset~q ),
	.datae(!\always5~0_combout ),
	.dataf(!\clear_crc~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~1 .extended_lut = "off";
defparam \always5~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \always5~1 .shared_arith = "off";

cyclonev_lcell_comb \enable_crc_calculation~0 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[2]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[1]~q ),
	.dataf(!\bit_counter|auto_generated|counter_reg_bit[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_crc_calculation~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_crc_calculation~0 .extended_lut = "off";
defparam \enable_crc_calculation~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \enable_crc_calculation~0 .shared_arith = "off";

cyclonev_lcell_comb \always5~2 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datab(!\enable_crc_storage~1_combout ),
	.datac(!\device_dclk_en_without_sdr~2_combout ),
	.datad(!\always5~0_combout ),
	.datae(!\enable_crc_calculation~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~2 .extended_lut = "off";
defparam \always5~2 .lut_mask = 64'hFF69FF96FF69FF96;
defparam \always5~2 .shared_arith = "off";

cyclonev_lcell_comb \enable_crc_storage~2 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\device_dclk_en_without_sdr~0_combout ),
	.datac(!\always5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_crc_storage~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_crc_storage~2 .extended_lut = "off";
defparam \enable_crc_storage~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \enable_crc_storage~2 .shared_arith = "off";

cyclonev_lcell_comb \enable_crc_change~0 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[2]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[1]~q ),
	.dataf(!\bit_counter|auto_generated|counter_reg_bit[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_crc_change~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_crc_change~0 .extended_lut = "off";
defparam \enable_crc_change~0 .lut_mask = 64'h6996966996696996;
defparam \enable_crc_change~0 .shared_arith = "off";

cyclonev_lcell_comb \crc_reg[14]~0 (
	.dataa(!\enable_crc_storage~2_combout ),
	.datab(!\always5~2_combout ),
	.datac(!\enable_crc_change~0_combout ),
	.datad(!\always5~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_reg[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_reg[14]~0 .extended_lut = "off";
defparam \crc_reg[14]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \crc_reg[14]~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~14 (
	.dataa(!irf_reg_0_1),
	.datab(!\Equal6~1_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal23~0_combout ),
	.datae(!\sdr~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~14 .extended_lut = "off";
defparam \comb~14 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \comb~14 .shared_arith = "off";

cyclonev_lcell_comb \comb~15 (
	.dataa(!irf_reg_0_1),
	.datab(!\Equal6~1_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal23~0_combout ),
	.datae(!\sdr~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~15 .extended_lut = "off";
defparam \comb~15 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \comb~15 .shared_arith = "off";

cyclonev_lcell_comb \comb~16 (
	.dataa(!\Equal1~0_combout ),
	.datab(!irf_reg_9_1),
	.datac(!irf_reg_11_1),
	.datad(!\Equal17~0_combout ),
	.datae(!\sdr~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~16 .extended_lut = "off";
defparam \comb~16 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \comb~16 .shared_arith = "off";

cyclonev_lcell_comb \crc_reg~1 (
	.dataa(!\enable_crc_storage~2_combout ),
	.datab(!\crc_reg[15]~q ),
	.datac(!\always5~2_combout ),
	.datad(!\enable_crc_change~0_combout ),
	.datae(!\always5~1_combout ),
	.dataf(!\crc_reg[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_reg~1 .extended_lut = "off";
defparam \crc_reg~1 .lut_mask = 64'hBFFFB3FFFFFFFFFF;
defparam \crc_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \crc_wire[12] (
	.dataa(!data1out_int),
	.datab(!\crc_reg[15]~q ),
	.datac(!\crc_reg[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_wire[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_wire[12] .extended_lut = "off";
defparam \crc_wire[12] .lut_mask = 64'h9696969696969696;
defparam \crc_wire[12] .shared_arith = "off";

cyclonev_lcell_comb \crc_wire[5] (
	.dataa(!data1out_int),
	.datab(!\crc_reg[15]~q ),
	.datac(!\crc_reg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_wire[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_wire[5] .extended_lut = "off";
defparam \crc_wire[5] .lut_mask = 64'h9696969696969696;
defparam \crc_wire[5] .shared_arith = "off";

cyclonev_lcell_comb \Equal26~1 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal26),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~1 .extended_lut = "off";
defparam \Equal26~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal26~1 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~15 (
	.dataa(!\adapted_tdo~5_combout ),
	.datab(!\adapted_tdo~6_combout ),
	.datac(!\adapted_tdo~10_combout ),
	.datad(!\adapted_tdo~13_combout ),
	.datae(!\adapted_tdo~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(adapted_tdo),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~15 .extended_lut = "off";
defparam \adapted_tdo~15 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \adapted_tdo~15 .shared_arith = "off";

dffeas single_scein(
	.clk(!altera_internal_jtag),
	.d(\device_dclk_en_without_sdr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(single_scein1),
	.prn(vcc));
defparam single_scein.is_wysiwyg = "true";
defparam single_scein.power_up = "low";

dffeas \sdoin~reg0 (
	.clk(!altera_internal_jtag),
	.d(\sdoin_wire~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sdoin),
	.prn(vcc));
defparam \sdoin~reg0 .is_wysiwyg = "true";
defparam \sdoin~reg0 .power_up = "low";

cyclonev_lcell_comb \data1in~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_io1_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(data1in),
	.sumout(),
	.cout(),
	.shareout());
defparam \data1in~0 .extended_lut = "off";
defparam \data1in~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \data1in~0 .shared_arith = "off";

cyclonev_lcell_comb \data2in~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_io2_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(data2in),
	.sumout(),
	.cout(),
	.shareout());
defparam \data2in~0 .extended_lut = "off";
defparam \data2in~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \data2in~0 .shared_arith = "off";

cyclonev_lcell_comb \data3in~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_io3_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(data3in),
	.sumout(),
	.cout(),
	.shareout());
defparam \data3in~0 .extended_lut = "off";
defparam \data3in~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \data3in~0 .shared_arith = "off";

cyclonev_lcell_comb \dclkin~0 (
	.dataa(!\device_dclk_en_reg~q ),
	.datab(!\dclkin_without_sdr~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dclkin),
	.sumout(),
	.cout(),
	.shareout());
defparam \dclkin~0 .extended_lut = "off";
defparam \dclkin~0 .lut_mask = 64'h7777777777777777;
defparam \dclkin~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal11~1 (
	.dataa(!irf_reg_1_1),
	.datab(!irf_reg_8_1),
	.datac(!irf_reg_10_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~1 .extended_lut = "off";
defparam \Equal11~1 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Equal11~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~2 (
	.dataa(!irf_reg_2_1),
	.datab(!irf_reg_7_1),
	.datac(!irf_reg_6_1),
	.datad(!irf_reg_3_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~2 .extended_lut = "off";
defparam \Equal5~2 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \Equal5~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal26~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_4_1),
	.datac(!irf_reg_5_1),
	.datad(!irf_reg_9_1),
	.datae(!irf_reg_11_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~0 .extended_lut = "off";
defparam \Equal26~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \Equal26~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_2_1),
	.datac(!irf_reg_7_1),
	.datad(!irf_reg_6_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~0 .extended_lut = "off";
defparam \Equal17~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal17~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal11~0 (
	.dataa(!irf_reg_4_1),
	.datab(!irf_reg_3_1),
	.datac(!irf_reg_5_1),
	.datad(!irf_reg_9_1),
	.datae(!irf_reg_11_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~0 .extended_lut = "off";
defparam \Equal11~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!irf_reg_1_1),
	.datab(!irf_reg_8_1),
	.datac(!irf_reg_10_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~0 (
	.dataa(!\Equal17~0_combout ),
	.datab(!\Equal11~0_combout ),
	.datac(!\Equal6~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal14~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!irf_reg_1_1),
	.datab(!irf_reg_4_1),
	.datac(!irf_reg_8_1),
	.datad(!irf_reg_10_1),
	.datae(!irf_reg_3_1),
	.dataf(!irf_reg_5_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!irf_reg_6_1),
	.datab(!irf_reg_9_1),
	.datac(!irf_reg_11_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal10~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_2_1),
	.datac(!irf_reg_7_1),
	.datad(!\Equal1~0_combout ),
	.datae(!\Equal1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal10~0 .extended_lut = "off";
defparam \Equal10~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \Equal10~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~1 (
	.dataa(!irf_reg_2_1),
	.datab(!irf_reg_7_1),
	.datac(!irf_reg_6_1),
	.datad(!irf_reg_9_1),
	.datae(!irf_reg_11_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~1 .extended_lut = "off";
defparam \Equal6~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal6~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!irf_reg_8_1),
	.datab(!irf_reg_10_1),
	.datac(!irf_reg_5_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_4_1),
	.datac(!irf_reg_3_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Equal16~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~1 (
	.dataa(!irf_reg_1_1),
	.datab(!\Equal6~1_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal16~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~1 .extended_lut = "off";
defparam \Equal16~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Equal16~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~0 (
	.dataa(!irf_reg_1_1),
	.datab(!irf_reg_8_1),
	.datac(!irf_reg_10_1),
	.datad(!\Equal17~0_combout ),
	.datae(!\Equal11~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~0 .extended_lut = "off";
defparam \Equal15~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \Equal15~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal11~2 (
	.dataa(!\Equal17~0_combout ),
	.datab(!\Equal11~0_combout ),
	.datac(!\Equal11~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~2 .extended_lut = "off";
defparam \Equal11~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal11~2 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~0 (
	.dataa(gnd),
	.datab(!\Equal10~0_combout ),
	.datac(!\Equal16~1_combout ),
	.datad(!\Equal15~0_combout ),
	.datae(!\Equal11~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~0 .extended_lut = "off";
defparam \adapted_tdo~0 .lut_mask = 64'hFFFFFFFCFFFFFFFC;
defparam \adapted_tdo~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~1 (
	.dataa(!irf_reg_4_1),
	.datab(!irf_reg_3_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~1 .extended_lut = "off";
defparam \Equal3~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~2 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_1_1),
	.datac(!\Equal6~1_combout ),
	.datad(!\Equal3~0_combout ),
	.datae(!\Equal3~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~2 .extended_lut = "off";
defparam \Equal3~2 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \Equal3~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!irf_reg_9_1),
	.datab(!irf_reg_11_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~1 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_2_1),
	.datac(!irf_reg_7_1),
	.datad(!irf_reg_6_1),
	.datae(!\Equal1~0_combout ),
	.dataf(!\Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~1 .extended_lut = "off";
defparam \adapted_tdo~1 .lut_mask = 64'hF7FDFFFFFFFFFFFF;
defparam \adapted_tdo~1 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~2 (
	.dataa(!\Equal3~2_combout ),
	.datab(!\adapted_tdo~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~2 .extended_lut = "off";
defparam \adapted_tdo~2 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \adapted_tdo~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~1 (
	.dataa(!irf_reg_1_1),
	.datab(!irf_reg_4_1),
	.datac(!irf_reg_8_1),
	.datad(!irf_reg_10_1),
	.datae(!irf_reg_9_1),
	.dataf(!irf_reg_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~1 .extended_lut = "off";
defparam \Equal5~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal5~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~3 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_5_1),
	.datac(!\Equal5~1_combout ),
	.datad(!\Equal5~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~3 .extended_lut = "off";
defparam \Equal5~3 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \Equal5~3 .shared_arith = "off";

dffeas bypass_out(
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bypass_out~q ),
	.prn(vcc));
defparam bypass_out.is_wysiwyg = "true";
defparam bypass_out.power_up = "low";

cyclonev_lcell_comb \Equal6~2 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_4_1),
	.datac(!irf_reg_3_1),
	.datad(!irf_reg_5_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~2 .extended_lut = "off";
defparam \Equal6~2 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \Equal6~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~3 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~0_combout ),
	.datac(!\Equal6~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~3 .extended_lut = "off";
defparam \Equal6~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal6~3 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~3 (
	.dataa(!\Equal5~3_combout ),
	.datab(!\powerful_reg|dffs[0]~q ),
	.datac(!Equal26),
	.datad(!\bypass_out~q ),
	.datae(!\Equal6~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~3 .extended_lut = "off";
defparam \adapted_tdo~3 .lut_mask = 64'hBFFFB3FFBFFFB3FF;
defparam \adapted_tdo~3 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~4 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\crc_shifter|dffs[0]~q ),
	.datac(!\Equal5~3_combout ),
	.datad(!\Equal6~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~4 .extended_lut = "off";
defparam \adapted_tdo~4 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \adapted_tdo~4 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~5 (
	.dataa(!\Equal14~0_combout ),
	.datab(!\adapted_tdo~0_combout ),
	.datac(!\adapted_tdo~2_combout ),
	.datad(!\adapted_tdo~3_combout ),
	.datae(!\adapted_tdo~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~5 .extended_lut = "off";
defparam \adapted_tdo~5 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \adapted_tdo~5 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~6 (
	.dataa(!\Equal14~0_combout ),
	.datab(!\adapted_tdo~0_combout ),
	.datac(!\data_speed_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.datad(!\adapted_tdo~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~6 .extended_lut = "off";
defparam \adapted_tdo~6 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \adapted_tdo~6 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~7 (
	.dataa(!\Equal10~0_combout ),
	.datab(!\Equal16~1_combout ),
	.datac(!\opcode_reg|dffs[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~7 .extended_lut = "off";
defparam \adapted_tdo~7 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \adapted_tdo~7 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~8 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\Equal10~0_combout ),
	.datac(!\Equal16~1_combout ),
	.datad(!\Equal15~0_combout ),
	.datae(!\Equal11~2_combout ),
	.dataf(!\rsiid_reg|dffs[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~8 .extended_lut = "off";
defparam \adapted_tdo~8 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \adapted_tdo~8 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~9 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\Equal10~0_combout ),
	.datac(!\Equal16~1_combout ),
	.datad(!\Equal15~0_combout ),
	.datae(!\Equal11~2_combout ),
	.dataf(!\rdi_reg|dffs[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~9 .extended_lut = "off";
defparam \adapted_tdo~9 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \adapted_tdo~9 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~10 (
	.dataa(!\adapted_tdo~7_combout ),
	.datab(!\rstatus_reg|dffs[0]~q ),
	.datac(!\Equal14~0_combout ),
	.datad(!\adapted_tdo~0_combout ),
	.datae(!\adapted_tdo~8_combout ),
	.dataf(!\adapted_tdo~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~10 .extended_lut = "off";
defparam \adapted_tdo~10 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \adapted_tdo~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal21~0 (
	.dataa(!\Equal1~0_combout ),
	.datab(!irf_reg_9_1),
	.datac(!irf_reg_11_1),
	.datad(!\Equal17~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~0 .extended_lut = "off";
defparam \Equal21~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \Equal21~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~1 (
	.dataa(!irf_reg_3_1),
	.datab(!irf_reg_5_1),
	.datac(!\Equal17~0_combout ),
	.datad(!\Equal5~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~1 .extended_lut = "off";
defparam \Equal17~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Equal17~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!irf_reg_2_1),
	.datab(!irf_reg_7_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!irf_reg_0_1),
	.datab(!\Equal1~0_combout ),
	.datac(!\Equal1~1_combout ),
	.datad(!\Equal4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal19~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\Equal1~0_combout ),
	.datac(!\Equal1~1_combout ),
	.datad(!\Equal4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal19~0 .extended_lut = "off";
defparam \Equal19~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Equal19~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~4 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_4_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~4 .extended_lut = "off";
defparam \Equal6~4 .lut_mask = 64'h7777777777777777;
defparam \Equal6~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal23~0 (
	.dataa(!irf_reg_1_1),
	.datab(!irf_reg_3_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~0 .extended_lut = "off";
defparam \Equal23~0 .lut_mask = 64'h7777777777777777;
defparam \Equal23~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal25~0 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~4_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal23~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal25~0 .extended_lut = "off";
defparam \Equal25~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal25~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal20~0 (
	.dataa(!irf_reg_9_1),
	.datab(!irf_reg_11_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~0 .extended_lut = "off";
defparam \Equal20~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Equal20~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal20~1 (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal17~0_combout ),
	.datac(!\Equal20~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~1 .extended_lut = "off";
defparam \Equal20~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal20~1 .shared_arith = "off";

cyclonev_lcell_comb \always8~0 (
	.dataa(!\Equal4~1_combout ),
	.datab(!\Equal19~0_combout ),
	.datac(!\Equal25~0_combout ),
	.datad(!\Equal20~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always8~0 .extended_lut = "off";
defparam \always8~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \always8~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal13~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_1_1),
	.datac(!\Equal6~1_combout ),
	.datad(!\Equal3~0_combout ),
	.datae(!\Equal3~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal13~0 .extended_lut = "off";
defparam \Equal13~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \Equal13~0 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~11 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_2_1),
	.datac(!irf_reg_7_1),
	.datad(!irf_reg_6_1),
	.datae(!\Equal1~0_combout ),
	.dataf(!\Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~11 .extended_lut = "off";
defparam \adapted_tdo~11 .lut_mask = 64'hFBFEFFFFFFFFFFFF;
defparam \adapted_tdo~11 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~12 (
	.dataa(!\Equal13~0_combout ),
	.datab(!\adapted_tdo~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~12 .extended_lut = "off";
defparam \adapted_tdo~12 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \adapted_tdo~12 .shared_arith = "off";

cyclonev_lcell_comb \adapted_tdo~13 (
	.dataa(gnd),
	.datab(!\Equal21~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(!\always8~0_combout ),
	.datae(!\adapted_tdo~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~13 .extended_lut = "off";
defparam \adapted_tdo~13 .lut_mask = 64'hFCFFFFFFFCFFFFFF;
defparam \adapted_tdo~13 .shared_arith = "off";

cyclonev_lcell_comb \push_rsiid_inst~0 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\Equal21~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\push_rsiid_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \push_rsiid_inst~0 .extended_lut = "off";
defparam \push_rsiid_inst~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \push_rsiid_inst~0 .shared_arith = "off";

cyclonev_lcell_comb \push_rdi_inst~0 (
	.dataa(!\Equal1~0_combout ),
	.datab(!irf_reg_9_1),
	.datac(!irf_reg_11_1),
	.datad(!\Equal17~0_combout ),
	.datae(!\en4b_reg|dffs[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\push_rdi_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \push_rdi_inst~0 .extended_lut = "off";
defparam \push_rdi_inst~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \push_rdi_inst~0 .shared_arith = "off";

cyclonev_lcell_comb sdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!state_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam sdr.extended_lut = "off";
defparam sdr.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam sdr.shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_2_1),
	.datac(!irf_reg_7_1),
	.datad(!irf_reg_6_1),
	.datae(!\Equal1~0_combout ),
	.dataf(!\Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \enable_crc_storage~1 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[10]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[9]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[8]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[7]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_crc_storage~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_crc_storage~1 .extended_lut = "off";
defparam \enable_crc_storage~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \enable_crc_storage~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan19~0 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datac(!\enable_crc_storage~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan19~0 .extended_lut = "off";
defparam \LessThan19~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \LessThan19~0 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~1 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_2_1),
	.datac(!irf_reg_7_1),
	.datad(!irf_reg_6_1),
	.datae(!\Equal1~0_combout ),
	.dataf(!\Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~1 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~1 .lut_mask = 64'hEFFEFFFFFFFFFFFF;
defparam \device_dclk_en_without_sdr~1 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~2 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~2 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~2 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \device_dclk_en_without_sdr~2 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~3 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datab(!\enable_crc_storage~1_combout ),
	.datac(!\device_dclk_en_without_sdr~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~3 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~3 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \device_dclk_en_without_sdr~3 .shared_arith = "off";

cyclonev_lcell_comb \enable_speed_write_data~0 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_speed_write_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_speed_write_data~0 .extended_lut = "off";
defparam \enable_speed_write_data~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \enable_speed_write_data~0 .shared_arith = "off";

cyclonev_lcell_comb \always4~0 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always4~0 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~4 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datac(!\enable_crc_storage~1_combout ),
	.datad(!\enable_speed_write_data~0_combout ),
	.datae(!\always4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~4 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~4 .lut_mask = 64'hBEFFFFFFBEFFFFFF;
defparam \device_dclk_en_without_sdr~4 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~5 (
	.dataa(!\Equal4~1_combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\LessThan19~0_combout ),
	.datad(!\device_dclk_en_without_sdr~1_combout ),
	.datae(!\device_dclk_en_without_sdr~3_combout ),
	.dataf(!\device_dclk_en_without_sdr~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~5 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~5 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \device_dclk_en_without_sdr~5 .shared_arith = "off";

cyclonev_lcell_comb \push_rsiid_inst~1 (
	.dataa(!\Equal1~0_combout ),
	.datab(!irf_reg_9_1),
	.datac(!irf_reg_11_1),
	.datad(!\Equal17~0_combout ),
	.datae(!\en4b_reg|dffs[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\push_rsiid_inst~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \push_rsiid_inst~1 .extended_lut = "off";
defparam \push_rsiid_inst~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \push_rsiid_inst~1 .shared_arith = "off";

cyclonev_lcell_comb \always4~1 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[10]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[9]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[8]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[7]~q ),
	.dataf(!\bit_counter|auto_generated|counter_reg_bit[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~1 .extended_lut = "off";
defparam \always4~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \always4~1 .shared_arith = "off";

cyclonev_lcell_comb \always4~2 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\always4~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~2 .extended_lut = "off";
defparam \always4~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always4~2 .shared_arith = "off";

cyclonev_lcell_comb \always4~3 (
	.dataa(!irf_reg_1_1),
	.datab(!\Equal6~1_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal16~0_combout ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.dataf(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~3 .extended_lut = "off";
defparam \always4~3 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \always4~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan20~0 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan20~0 .extended_lut = "off";
defparam \LessThan20~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \LessThan20~0 .shared_arith = "off";

cyclonev_lcell_comb \always4~4 (
	.dataa(!\LessThan20~0_combout ),
	.datab(!\always4~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~4 .extended_lut = "off";
defparam \always4~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always4~4 .shared_arith = "off";

cyclonev_lcell_comb \always4~5 (
	.dataa(!\Equal1~0_combout ),
	.datab(!\Equal17~0_combout ),
	.datac(!\Equal20~0_combout ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.dataf(!\always4~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~5 .extended_lut = "off";
defparam \always4~5 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \always4~5 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~6 (
	.dataa(!\push_rsiid_inst~1_combout ),
	.datab(!\Equal17~1_combout ),
	.datac(!\always4~2_combout ),
	.datad(!\always4~3_combout ),
	.datae(!\always4~4_combout ),
	.dataf(!\always4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~6 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~6 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \device_dclk_en_without_sdr~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal23~1 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_4_1),
	.datac(!\Equal6~1_combout ),
	.datad(!\Equal3~0_combout ),
	.datae(!\Equal23~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~1 .extended_lut = "off";
defparam \Equal23~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \Equal23~1 .shared_arith = "off";

cyclonev_lcell_comb \always4~6 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~4_combout ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal23~0_combout ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.dataf(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~6 .extended_lut = "off";
defparam \always4~6 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \always4~6 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~7 (
	.dataa(!\push_rdi_inst~0_combout ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datad(!\always4~1_combout ),
	.datae(!\Equal23~1_combout ),
	.dataf(!\always4~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~7 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~7 .lut_mask = 64'hFDFFF7FFF7FFFDFF;
defparam \device_dclk_en_without_sdr~7 .shared_arith = "off";

cyclonev_lcell_comb \data1out_reg~0 (
	.dataa(!\data1out_reg~q ),
	.datab(!\sdr~combout ),
	.datac(!data1out_int),
	.datad(!\device_dclk_en_without_sdr~5_combout ),
	.datae(!\device_dclk_en_without_sdr~6_combout ),
	.dataf(!\device_dclk_en_without_sdr~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data1out_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data1out_reg~0 .extended_lut = "off";
defparam \data1out_reg~0 .lut_mask = 64'h7FDFDF7FDF7F7FDF;
defparam \data1out_reg~0 .shared_arith = "off";

dffeas data1out_reg(
	.clk(altera_internal_jtag),
	.d(\data1out_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data1out_reg~q ),
	.prn(vcc));
defparam data1out_reg.is_wysiwyg = "true";
defparam data1out_reg.power_up = "low";

cyclonev_lcell_comb \adapted_tdo~14 (
	.dataa(!\push_rsiid_inst~0_combout ),
	.datab(!\push_rdi_inst~0_combout ),
	.datac(!\data1out_reg~q ),
	.datad(!\always8~0_combout ),
	.datae(!\data_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.dataf(!\adapted_tdo~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\adapted_tdo~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \adapted_tdo~14 .extended_lut = "off";
defparam \adapted_tdo~14 .lut_mask = 64'hFFFFFFFF9F6FFFFF;
defparam \adapted_tdo~14 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~8 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datad(!\enable_crc_storage~1_combout ),
	.datae(!\enable_speed_write_data~0_combout ),
	.dataf(!\always4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~8 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~8 .lut_mask = 64'hFFFFFFFFFFFF7FF7;
defparam \device_dclk_en_without_sdr~8 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~9 (
	.dataa(!\Equal4~1_combout ),
	.datab(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[11]~q ),
	.datad(!\enable_crc_storage~1_combout ),
	.datae(!\device_dclk_en_without_sdr~1_combout ),
	.dataf(!\device_dclk_en_without_sdr~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~9 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~9 .lut_mask = 64'hFFFFFFFFFDFFFFFF;
defparam \device_dclk_en_without_sdr~9 .shared_arith = "off";

cyclonev_lcell_comb \always4~7 (
	.dataa(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datab(!\always4~1_combout ),
	.datac(!\always4~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~7 .extended_lut = "off";
defparam \always4~7 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \always4~7 .shared_arith = "off";

cyclonev_lcell_comb \always4~8 (
	.dataa(!\push_rsiid_inst~1_combout ),
	.datab(!\Equal17~1_combout ),
	.datac(!\LessThan20~0_combout ),
	.datad(!\always4~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~8 .extended_lut = "off";
defparam \always4~8 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \always4~8 .shared_arith = "off";

cyclonev_lcell_comb \device_dclk_en_without_sdr~10 (
	.dataa(!\device_dclk_en_without_sdr~8_combout ),
	.datab(!\device_dclk_en_without_sdr~9_combout ),
	.datac(!\always4~7_combout ),
	.datad(!\always4~8_combout ),
	.datae(!\always4~5_combout ),
	.dataf(!\device_dclk_en_without_sdr~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~10 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~10 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \device_dclk_en_without_sdr~10 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~0 (
	.dataa(!\en4b_reg|dffs[0]~q ),
	.datab(!\Equal21~0_combout ),
	.datac(!\Equal16~1_combout ),
	.datad(!\opcode_reg|dffs[0]~q ),
	.datae(!\rdi_reg|dffs[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~0 .extended_lut = "off";
defparam \sdoin_wire~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sdoin_wire~0 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~1 (
	.dataa(!\push_rsiid_inst~0_combout ),
	.datab(!Equal26),
	.datac(!\device_dclk_en_without_sdr~1_combout ),
	.datad(!\sdoin_wire~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~1 .extended_lut = "off";
defparam \sdoin_wire~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \sdoin_wire~1 .shared_arith = "off";

cyclonev_lcell_comb \powerful_io0_reg~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_reg|dffs[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_io0_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \powerful_io0_reg~0 .extended_lut = "off";
defparam \powerful_io0_reg~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \powerful_io0_reg~0 .shared_arith = "off";

cyclonev_lcell_comb udr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!state_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\udr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam udr.extended_lut = "off";
defparam udr.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam udr.shared_arith = "off";

cyclonev_lcell_comb \powerful_ncs_reg~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\udr~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_ncs_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \powerful_ncs_reg~0 .extended_lut = "off";
defparam \powerful_ncs_reg~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \powerful_ncs_reg~0 .shared_arith = "off";

dffeas powerful_io0_reg(
	.clk(altera_internal_jtag),
	.d(\powerful_io0_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\powerful_ncs_reg~0_combout ),
	.q(\powerful_io0_reg~q ),
	.prn(vcc));
defparam powerful_io0_reg.is_wysiwyg = "true";
defparam powerful_io0_reg.power_up = "low";

cyclonev_lcell_comb \sdoin_wire~3 (
	.dataa(!\push_rsiid_inst~0_combout ),
	.datab(!\rsiid_reg|dffs[0]~q ),
	.datac(!Equal26),
	.datad(!\data_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.datae(!\device_dclk_en_without_sdr~1_combout ),
	.dataf(!\powerful_io0_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~3 .extended_lut = "off";
defparam \sdoin_wire~3 .lut_mask = 64'hBFFFFBFFFFFFFFFF;
defparam \sdoin_wire~3 .shared_arith = "off";

cyclonev_lcell_comb \comb~10 (
	.dataa(gnd),
	.datab(!\Equal21~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(!\Equal16~1_combout ),
	.datae(!\device_dclk_en_without_sdr~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~10 .extended_lut = "off";
defparam \comb~10 .lut_mask = 64'hFFFFFFFCFFFFFFFC;
defparam \comb~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal27~0 (
	.dataa(!\Equal1~0_combout ),
	.datab(!irf_reg_9_1),
	.datac(!irf_reg_11_1),
	.datad(!\Equal17~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal27~0 .extended_lut = "off";
defparam \Equal27~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal27~0 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~2 (
	.dataa(!\Equal25~0_combout ),
	.datab(!\aai_data_reg|dffs[0]~q ),
	.datac(!\ncso_reg|dffs[0]~q ),
	.datad(!\Equal27~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~2 .extended_lut = "off";
defparam \sdoin_wire~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sdoin_wire~2 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~6 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal4~1_combout ),
	.datac(!\aai_write_reg|dffs[0]~q ),
	.datad(!\rstatus_reg|dffs[0]~q ),
	.datae(!\Equal23~1_combout ),
	.dataf(!\Equal20~1_combout ),
	.datag(!\sdoin_wire~2_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~6 .extended_lut = "on";
defparam \sdoin_wire~6 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sdoin_wire~6 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~10 (
	.dataa(!\aai_write_reg|dffs[0]~q ),
	.datab(!\Equal23~1_combout ),
	.datac(!\sdoin_wire~2_combout ),
	.datad(!\Equal2~0_combout ),
	.datae(!\Equal4~1_combout ),
	.dataf(!\Equal20~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~10 .extended_lut = "off";
defparam \sdoin_wire~10 .lut_mask = 64'hDFFFFFFF1FFFFFFF;
defparam \sdoin_wire~10 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~5 (
	.dataa(!\data_speed_reg|dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.datab(!\sdoin_wire~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~5 .extended_lut = "off";
defparam \sdoin_wire~5 .lut_mask = 64'h7777777777777777;
defparam \sdoin_wire~5 .shared_arith = "off";

cyclonev_lcell_comb \sdoin_wire~4 (
	.dataa(!\sdoin_wire~1_combout ),
	.datab(!\sdoin_wire~3_combout ),
	.datac(!Equal26),
	.datad(!\comb~10_combout ),
	.datae(!\sdoin_wire~6_combout ),
	.dataf(!\sdoin_wire~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdoin_wire~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdoin_wire~4 .extended_lut = "off";
defparam \sdoin_wire~4 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \sdoin_wire~4 .shared_arith = "off";

cyclonev_lcell_comb \powerful_io1_reg~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_reg|dffs[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_io1_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \powerful_io1_reg~0 .extended_lut = "off";
defparam \powerful_io1_reg~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \powerful_io1_reg~0 .shared_arith = "off";

dffeas powerful_io1_reg(
	.clk(altera_internal_jtag),
	.d(\powerful_io1_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\powerful_ncs_reg~0_combout ),
	.q(\powerful_io1_reg~q ),
	.prn(vcc));
defparam powerful_io1_reg.is_wysiwyg = "true";
defparam powerful_io1_reg.power_up = "low";

cyclonev_lcell_comb \powerful_io2_reg~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_reg|dffs[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_io2_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \powerful_io2_reg~0 .extended_lut = "off";
defparam \powerful_io2_reg~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \powerful_io2_reg~0 .shared_arith = "off";

dffeas powerful_io2_reg(
	.clk(altera_internal_jtag),
	.d(\powerful_io2_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\powerful_ncs_reg~0_combout ),
	.q(\powerful_io2_reg~q ),
	.prn(vcc));
defparam powerful_io2_reg.is_wysiwyg = "true";
defparam powerful_io2_reg.power_up = "low";

cyclonev_lcell_comb \powerful_io3_reg~0 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\powerful_reg|dffs[0]~q ),
	.datad(!\Equal26~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_io3_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \powerful_io3_reg~0 .extended_lut = "off";
defparam \powerful_io3_reg~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \powerful_io3_reg~0 .shared_arith = "off";

dffeas powerful_io3_reg(
	.clk(altera_internal_jtag),
	.d(\powerful_io3_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\powerful_ncs_reg~0_combout ),
	.q(\powerful_io3_reg~q ),
	.prn(vcc));
defparam powerful_io3_reg.is_wysiwyg = "true";
defparam powerful_io3_reg.power_up = "low";

cyclonev_lcell_comb \device_dclk_en_without_sdr~11 (
	.dataa(!\push_rsiid_inst~0_combout ),
	.datab(!\Equal20~1_combout ),
	.datac(!\bit_counter|auto_generated|counter_reg_bit[5]~q ),
	.datad(!\bit_counter|auto_generated|counter_reg_bit[4]~q ),
	.datae(!\bit_counter|auto_generated|counter_reg_bit[3]~q ),
	.dataf(!\always4~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en_without_sdr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \device_dclk_en_without_sdr~11 .extended_lut = "off";
defparam \device_dclk_en_without_sdr~11 .lut_mask = 64'hFFFFFFFBFFFFFFFF;
defparam \device_dclk_en_without_sdr~11 .shared_arith = "off";

cyclonev_lcell_comb device_dclk_en(
	.dataa(!\sdr~combout ),
	.datab(!\device_dclk_en_without_sdr~8_combout ),
	.datac(!\device_dclk_en_without_sdr~9_combout ),
	.datad(!\always4~7_combout ),
	.datae(!\device_dclk_en_without_sdr~11_combout ),
	.dataf(!\device_dclk_en_without_sdr~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\device_dclk_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam device_dclk_en.extended_lut = "off";
defparam device_dclk_en.lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam device_dclk_en.shared_arith = "off";

dffeas device_dclk_en_reg(
	.clk(!altera_internal_jtag),
	.d(\device_dclk_en~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\device_dclk_en_reg~q ),
	.prn(vcc));
defparam device_dclk_en_reg.is_wysiwyg = "true";
defparam device_dclk_en_reg.power_up = "low";

cyclonev_lcell_comb \powerful_ncs_reg~1 (
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!\powerful_reg|dffs[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_ncs_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \powerful_ncs_reg~1 .extended_lut = "off";
defparam \powerful_ncs_reg~1 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \powerful_ncs_reg~1 .shared_arith = "off";

dffeas powerful_ncs_reg(
	.clk(altera_internal_jtag),
	.d(\powerful_ncs_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\powerful_ncs_reg~0_combout ),
	.q(\powerful_ncs_reg~q ),
	.prn(vcc));
defparam powerful_ncs_reg.is_wysiwyg = "true";
defparam powerful_ncs_reg.power_up = "low";

dffeas udr_reg(
	.clk(altera_internal_jtag),
	.d(\udr~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\udr_reg~q ),
	.prn(vcc));
defparam udr_reg.is_wysiwyg = "true";
defparam udr_reg.power_up = "low";

cyclonev_lcell_comb powerful_sck(
	.dataa(!\Equal11~1_combout ),
	.datab(!\Equal5~2_combout ),
	.datac(!\Equal26~0_combout ),
	.datad(!altera_internal_jtag),
	.datae(!\powerful_ncs_reg~q ),
	.dataf(!\udr_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\powerful_sck~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam powerful_sck.extended_lut = "off";
defparam powerful_sck.lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam powerful_sck.shared_arith = "off";

cyclonev_lcell_comb dclkin_without_sdr(
	.dataa(!altera_internal_jtag),
	.datab(!\powerful_sck~combout ),
	.datac(!Equal26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dclkin_without_sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam dclkin_without_sdr.extended_lut = "off";
defparam dclkin_without_sdr.lut_mask = 64'h5353535353535353;
defparam dclkin_without_sdr.shared_arith = "off";

endmodule

module SerialFlashLoader_lpm_counter_1 (
	counter_reg_bit_5,
	counter_reg_bit_11,
	counter_reg_bit_10,
	counter_reg_bit_9,
	counter_reg_bit_8,
	counter_reg_bit_7,
	counter_reg_bit_6,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	sdrs_reg,
	comb,
	counter_reg_bit_0,
	clock)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_5;
output 	counter_reg_bit_11;
output 	counter_reg_bit_10;
output 	counter_reg_bit_9;
output 	counter_reg_bit_8;
output 	counter_reg_bit_7;
output 	counter_reg_bit_6;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	sdrs_reg;
input 	comb;
output 	counter_reg_bit_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



SerialFlashLoader_cntr_88i auto_generated(
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_11(counter_reg_bit_11),
	.counter_reg_bit_10(counter_reg_bit_10),
	.counter_reg_bit_9(counter_reg_bit_9),
	.counter_reg_bit_8(counter_reg_bit_8),
	.counter_reg_bit_7(counter_reg_bit_7),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.sdrs_reg(sdrs_reg),
	.comb(comb),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock));

endmodule

module SerialFlashLoader_cntr_88i (
	counter_reg_bit_5,
	counter_reg_bit_11,
	counter_reg_bit_10,
	counter_reg_bit_9,
	counter_reg_bit_8,
	counter_reg_bit_7,
	counter_reg_bit_6,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	sdrs_reg,
	comb,
	counter_reg_bit_0,
	clock)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_5;
output 	counter_reg_bit_11;
output 	counter_reg_bit_10;
output 	counter_reg_bit_9;
output 	counter_reg_bit_8;
output 	counter_reg_bit_7;
output 	counter_reg_bit_6;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	sdrs_reg;
input 	comb;
output 	counter_reg_bit_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~COUT ;
wire \counter_comb_bita7~COUT ;
wire \counter_comb_bita8~COUT ;
wire \counter_comb_bita9~COUT ;
wire \counter_comb_bita10~COUT ;
wire \counter_comb_bita11~sumout ;
wire \counter_comb_bita10~sumout ;
wire \counter_comb_bita9~sumout ;
wire \counter_comb_bita8~sumout ;
wire \counter_comb_bita7~sumout ;
wire \counter_comb_bita6~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;


dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[11] (
	.clk(clock),
	.d(\counter_comb_bita11~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_11),
	.prn(vcc));
defparam \counter_reg_bit[11] .is_wysiwyg = "true";
defparam \counter_reg_bit[11] .power_up = "low";

dffeas \counter_reg_bit[10] (
	.clk(clock),
	.d(\counter_comb_bita10~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_10),
	.prn(vcc));
defparam \counter_reg_bit[10] .is_wysiwyg = "true";
defparam \counter_reg_bit[10] .power_up = "low";

dffeas \counter_reg_bit[9] (
	.clk(clock),
	.d(\counter_comb_bita9~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_9),
	.prn(vcc));
defparam \counter_reg_bit[9] .is_wysiwyg = "true";
defparam \counter_reg_bit[9] .power_up = "low";

dffeas \counter_reg_bit[8] (
	.clk(clock),
	.d(\counter_comb_bita8~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_8),
	.prn(vcc));
defparam \counter_reg_bit[8] .is_wysiwyg = "true";
defparam \counter_reg_bit[8] .power_up = "low";

dffeas \counter_reg_bit[7] (
	.clk(clock),
	.d(\counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_7),
	.prn(vcc));
defparam \counter_reg_bit[7] .is_wysiwyg = "true";
defparam \counter_reg_bit[7] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!sdrs_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(\counter_comb_bita5~COUT ),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita6(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita6~sumout ),
	.cout(\counter_comb_bita6~COUT ),
	.shareout());
defparam counter_comb_bita6.extended_lut = "off";
defparam counter_comb_bita6.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita6.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita7~sumout ),
	.cout(\counter_comb_bita7~COUT ),
	.shareout());
defparam counter_comb_bita7.extended_lut = "off";
defparam counter_comb_bita7.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita7.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita8(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita8~sumout ),
	.cout(\counter_comb_bita8~COUT ),
	.shareout());
defparam counter_comb_bita8.extended_lut = "off";
defparam counter_comb_bita8.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita8.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita9(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita9~sumout ),
	.cout(\counter_comb_bita9~COUT ),
	.shareout());
defparam counter_comb_bita9.extended_lut = "off";
defparam counter_comb_bita9.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita9.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita10(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita10~sumout ),
	.cout(\counter_comb_bita10~COUT ),
	.shareout());
defparam counter_comb_bita10.extended_lut = "off";
defparam counter_comb_bita10.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita10.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita11(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita11~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita11.extended_lut = "off";
defparam counter_comb_bita11.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita11.shared_arith = "off";

endmodule

module SerialFlashLoader_lpm_shiftreg_1 (
	reset,
	dffs_0,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	dffs_0;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs[23]~q ;
wire \dffs[22]~q ;
wire \dffs[21]~q ;
wire \dffs[20]~q ;
wire \dffs[19]~q ;
wire \dffs[18]~q ;
wire \dffs[17]~q ;
wire \dffs[16]~q ;
wire \dffs[15]~q ;
wire \dffs[14]~q ;
wire \dffs[13]~q ;
wire \dffs[12]~q ;
wire \dffs[11]~q ;
wire \dffs[10]~q ;
wire \dffs[9]~q ;
wire \dffs[8]~q ;
wire \dffs[7]~q ;
wire \dffs[6]~q ;
wire \dffs[5]~q ;
wire \dffs[4]~q ;
wire \dffs[3]~q ;
wire \dffs[2]~q ;
wire \dffs[1]~q ;


dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[23] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[23]~q ),
	.prn(vcc));
defparam \dffs[23] .is_wysiwyg = "true";
defparam \dffs[23] .power_up = "low";

dffeas \dffs[22] (
	.clk(clock),
	.d(\dffs[23]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[22]~q ),
	.prn(vcc));
defparam \dffs[22] .is_wysiwyg = "true";
defparam \dffs[22] .power_up = "low";

dffeas \dffs[21] (
	.clk(clock),
	.d(\dffs[22]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[21]~q ),
	.prn(vcc));
defparam \dffs[21] .is_wysiwyg = "true";
defparam \dffs[21] .power_up = "low";

dffeas \dffs[20] (
	.clk(clock),
	.d(\dffs[21]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[20]~q ),
	.prn(vcc));
defparam \dffs[20] .is_wysiwyg = "true";
defparam \dffs[20] .power_up = "low";

dffeas \dffs[19] (
	.clk(clock),
	.d(\dffs[20]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[19]~q ),
	.prn(vcc));
defparam \dffs[19] .is_wysiwyg = "true";
defparam \dffs[19] .power_up = "low";

dffeas \dffs[18] (
	.clk(clock),
	.d(\dffs[19]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[18]~q ),
	.prn(vcc));
defparam \dffs[18] .is_wysiwyg = "true";
defparam \dffs[18] .power_up = "low";

dffeas \dffs[17] (
	.clk(clock),
	.d(\dffs[18]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[17]~q ),
	.prn(vcc));
defparam \dffs[17] .is_wysiwyg = "true";
defparam \dffs[17] .power_up = "low";

dffeas \dffs[16] (
	.clk(clock),
	.d(\dffs[17]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[16]~q ),
	.prn(vcc));
defparam \dffs[16] .is_wysiwyg = "true";
defparam \dffs[16] .power_up = "low";

dffeas \dffs[15] (
	.clk(clock),
	.d(\dffs[16]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[15]~q ),
	.prn(vcc));
defparam \dffs[15] .is_wysiwyg = "true";
defparam \dffs[15] .power_up = "low";

dffeas \dffs[14] (
	.clk(clock),
	.d(\dffs[15]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[14]~q ),
	.prn(vcc));
defparam \dffs[14] .is_wysiwyg = "true";
defparam \dffs[14] .power_up = "low";

dffeas \dffs[13] (
	.clk(clock),
	.d(\dffs[14]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[13]~q ),
	.prn(vcc));
defparam \dffs[13] .is_wysiwyg = "true";
defparam \dffs[13] .power_up = "low";

dffeas \dffs[12] (
	.clk(clock),
	.d(\dffs[13]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[12]~q ),
	.prn(vcc));
defparam \dffs[12] .is_wysiwyg = "true";
defparam \dffs[12] .power_up = "low";

dffeas \dffs[11] (
	.clk(clock),
	.d(\dffs[12]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[11]~q ),
	.prn(vcc));
defparam \dffs[11] .is_wysiwyg = "true";
defparam \dffs[11] .power_up = "low";

dffeas \dffs[10] (
	.clk(clock),
	.d(\dffs[11]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[10]~q ),
	.prn(vcc));
defparam \dffs[10] .is_wysiwyg = "true";
defparam \dffs[10] .power_up = "low";

dffeas \dffs[9] (
	.clk(clock),
	.d(\dffs[10]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[9]~q ),
	.prn(vcc));
defparam \dffs[9] .is_wysiwyg = "true";
defparam \dffs[9] .power_up = "low";

dffeas \dffs[8] (
	.clk(clock),
	.d(\dffs[9]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[8]~q ),
	.prn(vcc));
defparam \dffs[8] .is_wysiwyg = "true";
defparam \dffs[8] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(\dffs[8]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[7]~q ),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(\dffs[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[6]~q ),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(\dffs[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[5]~q ),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(\dffs[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[4]~q ),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(\dffs[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[3]~q ),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(\dffs[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2]~q ),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(\dffs[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[1]~q ),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_2 (
	reset,
	dffs_0,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	dffs_0;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs[47]~q ;
wire \dffs[46]~q ;
wire \dffs[45]~q ;
wire \dffs[44]~q ;
wire \dffs[43]~q ;
wire \dffs[42]~q ;
wire \dffs[41]~q ;
wire \dffs[40]~q ;
wire \dffs[39]~q ;
wire \dffs[38]~q ;
wire \dffs[37]~q ;
wire \dffs[36]~q ;
wire \dffs[35]~q ;
wire \dffs[34]~q ;
wire \dffs[33]~q ;
wire \dffs[32]~q ;
wire \dffs[31]~q ;
wire \dffs[30]~q ;
wire \dffs[29]~q ;
wire \dffs[28]~q ;
wire \dffs[27]~q ;
wire \dffs[26]~q ;
wire \dffs[25]~q ;
wire \dffs[24]~q ;
wire \dffs[23]~q ;
wire \dffs[22]~q ;
wire \dffs[21]~q ;
wire \dffs[20]~q ;
wire \dffs[19]~q ;
wire \dffs[18]~q ;
wire \dffs[17]~q ;
wire \dffs[16]~q ;
wire \dffs[15]~q ;
wire \dffs[14]~q ;
wire \dffs[13]~q ;
wire \dffs[12]~q ;
wire \dffs[11]~q ;
wire \dffs[10]~q ;
wire \dffs[9]~q ;
wire \dffs[8]~q ;
wire \dffs[7]~q ;
wire \dffs[6]~q ;
wire \dffs[5]~q ;
wire \dffs[4]~q ;
wire \dffs[3]~q ;
wire \dffs[2]~q ;
wire \dffs[1]~q ;


dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[47] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[47]~q ),
	.prn(vcc));
defparam \dffs[47] .is_wysiwyg = "true";
defparam \dffs[47] .power_up = "low";

dffeas \dffs[46] (
	.clk(clock),
	.d(\dffs[47]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[46]~q ),
	.prn(vcc));
defparam \dffs[46] .is_wysiwyg = "true";
defparam \dffs[46] .power_up = "low";

dffeas \dffs[45] (
	.clk(clock),
	.d(\dffs[46]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[45]~q ),
	.prn(vcc));
defparam \dffs[45] .is_wysiwyg = "true";
defparam \dffs[45] .power_up = "low";

dffeas \dffs[44] (
	.clk(clock),
	.d(\dffs[45]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[44]~q ),
	.prn(vcc));
defparam \dffs[44] .is_wysiwyg = "true";
defparam \dffs[44] .power_up = "low";

dffeas \dffs[43] (
	.clk(clock),
	.d(\dffs[44]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[43]~q ),
	.prn(vcc));
defparam \dffs[43] .is_wysiwyg = "true";
defparam \dffs[43] .power_up = "low";

dffeas \dffs[42] (
	.clk(clock),
	.d(\dffs[43]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[42]~q ),
	.prn(vcc));
defparam \dffs[42] .is_wysiwyg = "true";
defparam \dffs[42] .power_up = "low";

dffeas \dffs[41] (
	.clk(clock),
	.d(\dffs[42]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[41]~q ),
	.prn(vcc));
defparam \dffs[41] .is_wysiwyg = "true";
defparam \dffs[41] .power_up = "low";

dffeas \dffs[40] (
	.clk(clock),
	.d(\dffs[41]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[40]~q ),
	.prn(vcc));
defparam \dffs[40] .is_wysiwyg = "true";
defparam \dffs[40] .power_up = "low";

dffeas \dffs[39] (
	.clk(clock),
	.d(\dffs[40]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[39]~q ),
	.prn(vcc));
defparam \dffs[39] .is_wysiwyg = "true";
defparam \dffs[39] .power_up = "low";

dffeas \dffs[38] (
	.clk(clock),
	.d(\dffs[39]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[38]~q ),
	.prn(vcc));
defparam \dffs[38] .is_wysiwyg = "true";
defparam \dffs[38] .power_up = "low";

dffeas \dffs[37] (
	.clk(clock),
	.d(\dffs[38]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[37]~q ),
	.prn(vcc));
defparam \dffs[37] .is_wysiwyg = "true";
defparam \dffs[37] .power_up = "low";

dffeas \dffs[36] (
	.clk(clock),
	.d(\dffs[37]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[36]~q ),
	.prn(vcc));
defparam \dffs[36] .is_wysiwyg = "true";
defparam \dffs[36] .power_up = "low";

dffeas \dffs[35] (
	.clk(clock),
	.d(\dffs[36]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[35]~q ),
	.prn(vcc));
defparam \dffs[35] .is_wysiwyg = "true";
defparam \dffs[35] .power_up = "low";

dffeas \dffs[34] (
	.clk(clock),
	.d(\dffs[35]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[34]~q ),
	.prn(vcc));
defparam \dffs[34] .is_wysiwyg = "true";
defparam \dffs[34] .power_up = "low";

dffeas \dffs[33] (
	.clk(clock),
	.d(\dffs[34]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[33]~q ),
	.prn(vcc));
defparam \dffs[33] .is_wysiwyg = "true";
defparam \dffs[33] .power_up = "low";

dffeas \dffs[32] (
	.clk(clock),
	.d(\dffs[33]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[32]~q ),
	.prn(vcc));
defparam \dffs[32] .is_wysiwyg = "true";
defparam \dffs[32] .power_up = "low";

dffeas \dffs[31] (
	.clk(clock),
	.d(\dffs[32]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[31]~q ),
	.prn(vcc));
defparam \dffs[31] .is_wysiwyg = "true";
defparam \dffs[31] .power_up = "low";

dffeas \dffs[30] (
	.clk(clock),
	.d(\dffs[31]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[30]~q ),
	.prn(vcc));
defparam \dffs[30] .is_wysiwyg = "true";
defparam \dffs[30] .power_up = "low";

dffeas \dffs[29] (
	.clk(clock),
	.d(\dffs[30]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[29]~q ),
	.prn(vcc));
defparam \dffs[29] .is_wysiwyg = "true";
defparam \dffs[29] .power_up = "low";

dffeas \dffs[28] (
	.clk(clock),
	.d(\dffs[29]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[28]~q ),
	.prn(vcc));
defparam \dffs[28] .is_wysiwyg = "true";
defparam \dffs[28] .power_up = "low";

dffeas \dffs[27] (
	.clk(clock),
	.d(\dffs[28]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[27]~q ),
	.prn(vcc));
defparam \dffs[27] .is_wysiwyg = "true";
defparam \dffs[27] .power_up = "low";

dffeas \dffs[26] (
	.clk(clock),
	.d(\dffs[27]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[26]~q ),
	.prn(vcc));
defparam \dffs[26] .is_wysiwyg = "true";
defparam \dffs[26] .power_up = "low";

dffeas \dffs[25] (
	.clk(clock),
	.d(\dffs[26]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[25]~q ),
	.prn(vcc));
defparam \dffs[25] .is_wysiwyg = "true";
defparam \dffs[25] .power_up = "low";

dffeas \dffs[24] (
	.clk(clock),
	.d(\dffs[25]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[24]~q ),
	.prn(vcc));
defparam \dffs[24] .is_wysiwyg = "true";
defparam \dffs[24] .power_up = "low";

dffeas \dffs[23] (
	.clk(clock),
	.d(\dffs[24]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[23]~q ),
	.prn(vcc));
defparam \dffs[23] .is_wysiwyg = "true";
defparam \dffs[23] .power_up = "low";

dffeas \dffs[22] (
	.clk(clock),
	.d(\dffs[23]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[22]~q ),
	.prn(vcc));
defparam \dffs[22] .is_wysiwyg = "true";
defparam \dffs[22] .power_up = "low";

dffeas \dffs[21] (
	.clk(clock),
	.d(\dffs[22]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[21]~q ),
	.prn(vcc));
defparam \dffs[21] .is_wysiwyg = "true";
defparam \dffs[21] .power_up = "low";

dffeas \dffs[20] (
	.clk(clock),
	.d(\dffs[21]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[20]~q ),
	.prn(vcc));
defparam \dffs[20] .is_wysiwyg = "true";
defparam \dffs[20] .power_up = "low";

dffeas \dffs[19] (
	.clk(clock),
	.d(\dffs[20]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[19]~q ),
	.prn(vcc));
defparam \dffs[19] .is_wysiwyg = "true";
defparam \dffs[19] .power_up = "low";

dffeas \dffs[18] (
	.clk(clock),
	.d(\dffs[19]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[18]~q ),
	.prn(vcc));
defparam \dffs[18] .is_wysiwyg = "true";
defparam \dffs[18] .power_up = "low";

dffeas \dffs[17] (
	.clk(clock),
	.d(\dffs[18]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[17]~q ),
	.prn(vcc));
defparam \dffs[17] .is_wysiwyg = "true";
defparam \dffs[17] .power_up = "low";

dffeas \dffs[16] (
	.clk(clock),
	.d(\dffs[17]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[16]~q ),
	.prn(vcc));
defparam \dffs[16] .is_wysiwyg = "true";
defparam \dffs[16] .power_up = "low";

dffeas \dffs[15] (
	.clk(clock),
	.d(\dffs[16]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[15]~q ),
	.prn(vcc));
defparam \dffs[15] .is_wysiwyg = "true";
defparam \dffs[15] .power_up = "low";

dffeas \dffs[14] (
	.clk(clock),
	.d(\dffs[15]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[14]~q ),
	.prn(vcc));
defparam \dffs[14] .is_wysiwyg = "true";
defparam \dffs[14] .power_up = "low";

dffeas \dffs[13] (
	.clk(clock),
	.d(\dffs[14]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[13]~q ),
	.prn(vcc));
defparam \dffs[13] .is_wysiwyg = "true";
defparam \dffs[13] .power_up = "low";

dffeas \dffs[12] (
	.clk(clock),
	.d(\dffs[13]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[12]~q ),
	.prn(vcc));
defparam \dffs[12] .is_wysiwyg = "true";
defparam \dffs[12] .power_up = "low";

dffeas \dffs[11] (
	.clk(clock),
	.d(\dffs[12]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[11]~q ),
	.prn(vcc));
defparam \dffs[11] .is_wysiwyg = "true";
defparam \dffs[11] .power_up = "low";

dffeas \dffs[10] (
	.clk(clock),
	.d(\dffs[11]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[10]~q ),
	.prn(vcc));
defparam \dffs[10] .is_wysiwyg = "true";
defparam \dffs[10] .power_up = "low";

dffeas \dffs[9] (
	.clk(clock),
	.d(\dffs[10]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[9]~q ),
	.prn(vcc));
defparam \dffs[9] .is_wysiwyg = "true";
defparam \dffs[9] .power_up = "low";

dffeas \dffs[8] (
	.clk(clock),
	.d(\dffs[9]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[8]~q ),
	.prn(vcc));
defparam \dffs[8] .is_wysiwyg = "true";
defparam \dffs[8] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(\dffs[8]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[7]~q ),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(\dffs[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[6]~q ),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(\dffs[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[5]~q ),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(\dffs[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[4]~q ),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(\dffs[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[3]~q ),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(\dffs[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2]~q ),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(\dffs[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[1]~q ),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_3 (
	dffs_0,
	reset,
	counter_reg_bit_5,
	device_dclk_en_without_sdr,
	comb,
	enable_crc_storage,
	always5,
	enable,
	crc_shifter_input,
	clock)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
input 	reset;
input 	counter_reg_bit_5;
input 	device_dclk_en_without_sdr;
input 	comb;
input 	enable_crc_storage;
input 	always5;
input 	enable;
input 	crc_shifter_input;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1_sumout ;
wire \dffs_rtl_0|auto_generated|dffe7~0_combout ;
wire \dffs_rtl_0|auto_generated|dffe7~q ;
wire \dffs[8191]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1_sumout ;
wire \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ;
wire \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ;
wire \dffs_rtl_0|auto_generated|op_2~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \dffs_rtl_0|auto_generated|op_1~1_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[0]~q ;
wire \dffs_rtl_0|auto_generated|cmpr4_aeb_int~2_combout ;
wire \dffs_rtl_0|auto_generated|op_1~2 ;
wire \dffs_rtl_0|auto_generated|op_1~5_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~q ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \dffs_rtl_0|auto_generated|op_1~6 ;
wire \dffs_rtl_0|auto_generated|op_1~9_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[2]~q ;
wire \dffs_rtl_0|auto_generated|op_1~10 ;
wire \dffs_rtl_0|auto_generated|op_1~13_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[3]~q ;
wire \dffs_rtl_0|auto_generated|op_1~14 ;
wire \dffs_rtl_0|auto_generated|op_1~17_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[4]~q ;
wire \dffs_rtl_0|auto_generated|op_1~18 ;
wire \dffs_rtl_0|auto_generated|op_1~21_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[5]~q ;
wire \dffs_rtl_0|auto_generated|op_1~22 ;
wire \dffs_rtl_0|auto_generated|op_1~25_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[6]~q ;
wire \dffs_rtl_0|auto_generated|op_1~26 ;
wire \dffs_rtl_0|auto_generated|op_1~29_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[7]~q ;
wire \dffs_rtl_0|auto_generated|op_1~30 ;
wire \dffs_rtl_0|auto_generated|op_1~33_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[8]~q ;
wire \dffs_rtl_0|auto_generated|op_1~34 ;
wire \dffs_rtl_0|auto_generated|op_1~37_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[9]~q ;
wire \dffs_rtl_0|auto_generated|op_1~38 ;
wire \dffs_rtl_0|auto_generated|op_1~41_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[10]~q ;
wire \dffs_rtl_0|auto_generated|op_1~42 ;
wire \dffs_rtl_0|auto_generated|op_1~45_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[11]~q ;
wire \dffs_rtl_0|auto_generated|op_1~46 ;
wire \dffs_rtl_0|auto_generated|op_1~49_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[12]~q ;
wire \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ;

wire [143:0] \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ;

assign \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout  = \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus [0];

dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 (
	.dataa(!counter_reg_bit_5),
	.datab(!device_dclk_en_without_sdr),
	.datac(!comb),
	.datad(!enable_crc_storage),
	.datae(!always5),
	.dataf(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit12 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1 .lut_mask = 64'h0000000000000000;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe7~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita12~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe7~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe7~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe7 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|dffe7~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe7~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe7 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe7 .power_up = "low";

dffeas \dffs[8191] (
	.clk(clock),
	.d(crc_shifter_input),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[8191]~q ),
	.prn(vcc));
defparam \dffs[8191] .is_wysiwyg = "true";
defparam \dffs[8191] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1 .lut_mask = 64'h0000000000000000;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datad(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \dffs_rtl_0|auto_generated|op_2~0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita12~1_sumout ),
	.datad(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cmpr4_aeb_int~2 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cmpr4_aeb_int~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~2 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~2 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~5 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~2_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h000055FF000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\dffs_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\dffs_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~9 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~2_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~14 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~17_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~18 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~17 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~17 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[4]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[4] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~21_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~22 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~21 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~21 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[5]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[5] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~25_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~26 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~25 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~25 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[6]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[6] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~29_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~30 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~29 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~29 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[7]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[7] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~33_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~34 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~33 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~33 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~33 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[8]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[8] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~37_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~38 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~37 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~37 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~37 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[9]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[9] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~41_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~42 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~41 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~41 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~41 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[10]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[10] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~45_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~46 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~45 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~45 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~45 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[11]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[11] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~49_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~49 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~49 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~49 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[12] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[12]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[12] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[12] .power_up = "low";

cyclonev_ram_block \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock),
	.clk1(clock),
	.ena0(enable),
	.ena1(enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\dffs_rtl_0|auto_generated|dffe7~q ),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dffs[8191]~q }),
	.portaaddr({gnd,gnd,gnd,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[12]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,\dffs_rtl_0|auto_generated|dffe3a[12]~q ,\dffs_rtl_0|auto_generated|dffe3a[11]~q ,\dffs_rtl_0|auto_generated|dffe3a[10]~q ,\dffs_rtl_0|auto_generated|dffe3a[9]~q ,\dffs_rtl_0|auto_generated|dffe3a[8]~q ,\dffs_rtl_0|auto_generated|dffe3a[7]~q ,
\dffs_rtl_0|auto_generated|dffe3a[6]~q ,\dffs_rtl_0|auto_generated|dffe3a[5]~q ,\dffs_rtl_0|auto_generated|dffe3a[4]~q ,\dffs_rtl_0|auto_generated|dffe3a[3]~q ,\dffs_rtl_0|auto_generated|dffe3a[2]~q ,\dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,
\dffs_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_core_clock_enable = "ena0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_input_clock_enable = "ena0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk1_output_clock_enable = "ena1";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_offset_in_bits = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_width_in_bits = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .logical_ram_name = "altera_serial_flash_loader:serial_flash_loader_0|altserial_flash_loader:altserial_flash_loader_component|alt_sfl_enhanced:\\ENHANCED_PGM_QUAD:sfl_inst_enhanced|lpm_shiftreg:crc_shifter|altshift_taps:dffs_rtl_0|shift_taps_ka31:auto_generated|altsyncram_7pc1:altsyncram5|ALTSYNCRAM";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .mixed_port_feed_through_mode = "dont_care";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .operation_mode = "dual_port";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_width = 13;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clock = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_address = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_bit_number = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_last_address = 8189;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_depth = 8190;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clock = "clock0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_width = 13;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clear = "clear0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clock = "clock1";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_address = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_bit_number = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_last_address = 8189;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_depth = 8190;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_enable_clock = "clock0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .ram_block_type = "auto";

endmodule

module SerialFlashLoader_lpm_shiftreg_4 (
	ram_block8a0,
	Equal19,
	Equal13,
	adapted_tdo,
	sdr,
	reset,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	ram_block8a0;
input 	Equal19;
input 	Equal13;
input 	adapted_tdo;
input 	sdr;
input 	reset;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ;
wire \dffs_rtl_0|auto_generated|dffe7~0_combout ;
wire \dffs_rtl_0|auto_generated|dffe7~q ;
wire \dffs[2079]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1_sumout ;
wire \dffs_rtl_0|auto_generated|op_2~0_combout ;
wire \dffs_rtl_0|auto_generated|op_2~1_combout ;
wire \dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \dffs_rtl_0|auto_generated|op_2~2_combout ;
wire \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ;
wire \dffs_rtl_0|auto_generated|op_1~1_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[0]~q ;
wire \dffs_rtl_0|auto_generated|op_1~2 ;
wire \dffs_rtl_0|auto_generated|op_1~5_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~q ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \dffs_rtl_0|auto_generated|op_1~6 ;
wire \dffs_rtl_0|auto_generated|op_1~9_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[2]~q ;
wire \dffs_rtl_0|auto_generated|op_1~10 ;
wire \dffs_rtl_0|auto_generated|op_1~13_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[3]~q ;
wire \dffs_rtl_0|auto_generated|op_1~14 ;
wire \dffs_rtl_0|auto_generated|op_1~17_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[4]~q ;
wire \dffs_rtl_0|auto_generated|op_1~18 ;
wire \dffs_rtl_0|auto_generated|op_1~21_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[5]~q ;
wire \dffs_rtl_0|auto_generated|op_1~22 ;
wire \dffs_rtl_0|auto_generated|op_1~25_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[6]~q ;
wire \dffs_rtl_0|auto_generated|op_1~26 ;
wire \dffs_rtl_0|auto_generated|op_1~29_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[7]~q ;
wire \dffs_rtl_0|auto_generated|op_1~30 ;
wire \dffs_rtl_0|auto_generated|op_1~33_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[8]~q ;
wire \dffs_rtl_0|auto_generated|op_1~34 ;
wire \dffs_rtl_0|auto_generated|op_1~37_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[9]~q ;
wire \dffs_rtl_0|auto_generated|op_1~38 ;
wire \dffs_rtl_0|auto_generated|op_1~41_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[10]~q ;
wire \dffs_rtl_0|auto_generated|op_1~42 ;
wire \dffs_rtl_0|auto_generated|op_1~45_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[11]~q ;

wire [143:0] \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ;

assign ram_block8a0 = \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus [0];

cyclonev_ram_block \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock),
	.clk1(clock),
	.ena0(enable),
	.ena1(enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\dffs_rtl_0|auto_generated|dffe7~q ),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dffs[2079]~q }),
	.portaaddr({gnd,gnd,gnd,gnd,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,\dffs_rtl_0|auto_generated|dffe3a[11]~q ,\dffs_rtl_0|auto_generated|dffe3a[10]~q ,\dffs_rtl_0|auto_generated|dffe3a[9]~q ,\dffs_rtl_0|auto_generated|dffe3a[8]~q ,\dffs_rtl_0|auto_generated|dffe3a[7]~q ,\dffs_rtl_0|auto_generated|dffe3a[6]~q ,
\dffs_rtl_0|auto_generated|dffe3a[5]~q ,\dffs_rtl_0|auto_generated|dffe3a[4]~q ,\dffs_rtl_0|auto_generated|dffe3a[3]~q ,\dffs_rtl_0|auto_generated|dffe3a[2]~q ,\dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\dffs_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_core_clock_enable = "ena0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_input_clock_enable = "ena0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk1_output_clock_enable = "ena1";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_offset_in_bits = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_width_in_bits = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .logical_ram_name = "altera_serial_flash_loader:serial_flash_loader_0|altserial_flash_loader:altserial_flash_loader_component|alt_sfl_enhanced:\\ENHANCED_PGM_QUAD:sfl_inst_enhanced|lpm_shiftreg:data_reg|altshift_taps:dffs_rtl_0|shift_taps_la31:auto_generated|altsyncram_5pc1:altsyncram5|ALTSYNCRAM";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .mixed_port_feed_through_mode = "dont_care";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .operation_mode = "dual_port";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_width = 12;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clock = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_address = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_bit_number = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_last_address = 2078;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_depth = 2079;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clock = "clock0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_width = 12;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clear = "clear0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clock = "clock1";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_address = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_bit_number = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_last_address = 2078;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_depth = 2079;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_enable_clock = "clock0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .ram_block_type = "auto";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 (
	.dataa(!Equal19),
	.datab(!Equal13),
	.datac(!sdr),
	.datad(!adapted_tdo),
	.datae(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 .lut_mask = 64'h0000000000000000;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe7~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe7~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe7~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe7 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|dffe7~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe7~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe7 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe7 .power_up = "low";

dffeas \dffs[2079] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2079]~q ),
	.prn(vcc));
defparam \dffs[2079] .is_wysiwyg = "true";
defparam \dffs[2079] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 .lut_mask = 64'h0000000000000000;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.dataf(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \dffs_rtl_0|auto_generated|op_2~0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~1 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \dffs_rtl_0|auto_generated|op_2~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1_sumout ),
	.datae(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.dataf(!\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~2 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datad(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datae(!\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~2 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \dffs_rtl_0|auto_generated|op_2~2 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datad(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datae(!\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~1 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h000055FF000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~5 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h000055FF000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\dffs_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\dffs_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~9 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~14 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~17_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~18 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~17 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~17 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[4]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[4] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~21 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~21_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~22 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~21 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~21 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~21 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[5]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[5] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~25 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~25_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~26 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~25 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~25 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~25 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[6]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[6] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~29 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~29_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~30 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~29 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~29 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~29 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[7]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[7] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~33 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~33_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~34 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~33 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~33 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~33 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[8]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[8] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~37 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~37_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~38 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~37 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~37 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~37 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[9]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[9] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~41 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~41_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~42 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~41 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~41 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~41 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[10]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[10] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~45_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~45 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~45 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~45 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[11]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[11] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_5 (
	ram_block8a0,
	Equal3,
	adapted_tdo,
	Equal4,
	sdr,
	reset,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	ram_block8a0;
input 	Equal3;
input 	adapted_tdo;
input 	Equal4;
input 	sdr;
input 	reset;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ;
wire \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ;
wire \dffs_rtl_0|auto_generated|dffe7~0_combout ;
wire \dffs_rtl_0|auto_generated|dffe7~q ;
wire \dffs[2107]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1_sumout ;
wire \dffs_rtl_0|auto_generated|op_2~0_combout ;
wire \dffs_rtl_0|auto_generated|op_2~1_combout ;
wire \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ;
wire \dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \dffs_rtl_0|auto_generated|op_2~2_combout ;
wire \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ;
wire \dffs_rtl_0|auto_generated|op_1~1_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[0]~q ;
wire \dffs_rtl_0|auto_generated|op_1~2 ;
wire \dffs_rtl_0|auto_generated|op_1~5_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~q ;
wire \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \dffs_rtl_0|auto_generated|op_1~6 ;
wire \dffs_rtl_0|auto_generated|op_1~9_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[2]~q ;
wire \dffs_rtl_0|auto_generated|op_1~10 ;
wire \dffs_rtl_0|auto_generated|op_1~13_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[3]~q ;
wire \dffs_rtl_0|auto_generated|op_1~14 ;
wire \dffs_rtl_0|auto_generated|op_1~17_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[4]~q ;
wire \dffs_rtl_0|auto_generated|op_1~18 ;
wire \dffs_rtl_0|auto_generated|op_1~21_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[5]~q ;
wire \dffs_rtl_0|auto_generated|op_1~22 ;
wire \dffs_rtl_0|auto_generated|op_1~25_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[6]~q ;
wire \dffs_rtl_0|auto_generated|op_1~26 ;
wire \dffs_rtl_0|auto_generated|op_1~29_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[7]~q ;
wire \dffs_rtl_0|auto_generated|op_1~30 ;
wire \dffs_rtl_0|auto_generated|op_1~33_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[8]~q ;
wire \dffs_rtl_0|auto_generated|op_1~34 ;
wire \dffs_rtl_0|auto_generated|op_1~37_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[9]~q ;
wire \dffs_rtl_0|auto_generated|op_1~38 ;
wire \dffs_rtl_0|auto_generated|op_1~41_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[10]~q ;
wire \dffs_rtl_0|auto_generated|op_1~42 ;
wire \dffs_rtl_0|auto_generated|op_1~45_sumout ;
wire \dffs_rtl_0|auto_generated|dffe3a[11]~q ;

wire [143:0] \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ;

assign ram_block8a0 = \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus [0];

cyclonev_ram_block \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock),
	.clk1(clock),
	.ena0(enable),
	.ena1(enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\dffs_rtl_0|auto_generated|dffe7~q ),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dffs[2107]~q }),
	.portaaddr({gnd,gnd,gnd,gnd,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,
\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,\dffs_rtl_0|auto_generated|dffe3a[11]~q ,\dffs_rtl_0|auto_generated|dffe3a[10]~q ,\dffs_rtl_0|auto_generated|dffe3a[9]~q ,\dffs_rtl_0|auto_generated|dffe3a[8]~q ,\dffs_rtl_0|auto_generated|dffe3a[7]~q ,\dffs_rtl_0|auto_generated|dffe3a[6]~q ,
\dffs_rtl_0|auto_generated|dffe3a[5]~q ,\dffs_rtl_0|auto_generated|dffe3a[4]~q ,\dffs_rtl_0|auto_generated|dffe3a[3]~q ,\dffs_rtl_0|auto_generated|dffe3a[2]~q ,\dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\dffs_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_core_clock_enable = "ena0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_input_clock_enable = "ena0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk1_output_clock_enable = "ena1";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_offset_in_bits = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_width_in_bits = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .logical_ram_name = "altera_serial_flash_loader:serial_flash_loader_0|altserial_flash_loader:altserial_flash_loader_component|alt_sfl_enhanced:\\ENHANCED_PGM_QUAD:sfl_inst_enhanced|lpm_shiftreg:data_speed_reg|altshift_taps:dffs_rtl_0|shift_taps_ca31:auto_generated|altsyncram_loc1:altsyncram5|ALTSYNCRAM";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .mixed_port_feed_through_mode = "dont_care";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .operation_mode = "dual_port";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_width = 12;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clock = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_address = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_bit_number = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_last_address = 2106;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_depth = 2107;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clear = "none";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clock = "clock0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_width = 12;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clear = "clear0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clock = "clock1";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_address = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_bit_number = 0;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_last_address = 2106;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_depth = 2107;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_width = 1;
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_enable_clock = "clock0";
defparam \dffs_rtl_0|auto_generated|altsyncram5|ram_block8a0 .ram_block_type = "auto";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 (
	.dataa(!Equal4),
	.datab(!Equal3),
	.datac(!sdr),
	.datad(!adapted_tdo),
	.datae(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit1 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit2 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit3 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit4 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit5 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit6 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit7 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit8 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit9 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~sumout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit10 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .lut_mask = 64'h000000000000FF00;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_reg_bit11 .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 .lut_mask = 64'h0000000000000000;
defparam \dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe7~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr6|counter_comb_bita11~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe7~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe7~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe7 (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|dffe7~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe7~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe7 .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe7 .power_up = "low";

dffeas \dffs[2107] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2107]~q ),
	.prn(vcc));
defparam \dffs[2107] .is_wysiwyg = "true";
defparam \dffs[2107] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita7~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita8~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita9~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita10~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ),
	.cout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 .lut_mask = 64'h0000000000000000;
defparam \dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \dffs_rtl_0|auto_generated|op_2~0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~1 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \dffs_rtl_0|auto_generated|op_2~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~0 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita11~1_sumout ),
	.datac(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datad(!\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.datae(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \dffs_rtl_0|auto_generated|cntr1|cout_actual .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dffs_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_2~2 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.dataf(!\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_2~2 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_2~2 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \dffs_rtl_0|auto_generated|op_2~2 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 (
	.dataa(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(!\dffs_rtl_0|auto_generated|op_2~0_combout ),
	.datac(!\dffs_rtl_0|auto_generated|op_2~1_combout ),
	.datad(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \dffs_rtl_0|auto_generated|cmpr4_aeb_int~1 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~1 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h000055FF000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[0] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~5 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h000055FF000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\dffs_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[1] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\dffs_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffs_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[2] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~13 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~14 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[3] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~17_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~18 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~17 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~17 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[4] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[4]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[4] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~21_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~22 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~21 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~21 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[5] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[5]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[5] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[5] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~25 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[6]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~25_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~26 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~25 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~25 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~25 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[6] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[6]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[6] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[6] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~29 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[7]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~29_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~30 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~29 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~29 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~29 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[7] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[7]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[7] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[7] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~33 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[8]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~33_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~34 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~33 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~33 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~33 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[8] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[8]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[8] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[8] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~37 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[9]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~37_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~38 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~37 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~37 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~37 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[9] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[9]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[9] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[9] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~41 (
	.dataa(!\dffs_rtl_0|auto_generated|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[10]~q ),
	.datae(gnd),
	.dataf(!\dffs_rtl_0|auto_generated|cmpr4_aeb_int~1_combout ),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~41_sumout ),
	.cout(\dffs_rtl_0|auto_generated|op_1~42 ),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~41 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~41 .lut_mask = 64'h0000FFAA000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~41 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[10] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[10]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[10] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[10] .power_up = "low";

cyclonev_lcell_comb \dffs_rtl_0|auto_generated|op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dffs_rtl_0|auto_generated|cntr1|counter_reg_bit[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dffs_rtl_0|auto_generated|op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dffs_rtl_0|auto_generated|op_1~45_sumout ),
	.cout(),
	.shareout());
defparam \dffs_rtl_0|auto_generated|op_1~45 .extended_lut = "off";
defparam \dffs_rtl_0|auto_generated|op_1~45 .lut_mask = 64'h00000000000000FF;
defparam \dffs_rtl_0|auto_generated|op_1~45 .shared_arith = "off";

dffeas \dffs_rtl_0|auto_generated|dffe3a[11] (
	.clk(clock),
	.d(\dffs_rtl_0|auto_generated|op_1~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs_rtl_0|auto_generated|dffe3a[11]~q ),
	.prn(vcc));
defparam \dffs_rtl_0|auto_generated|dffe3a[11] .is_wysiwyg = "true";
defparam \dffs_rtl_0|auto_generated|dffe3a[11] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_6 (
	dffs_0,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffs[0] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_7 (
	dffs_0,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs[7]~q ;
wire \dffs[6]~q ;
wire \dffs[5]~q ;
wire \dffs[4]~q ;
wire \dffs[3]~q ;
wire \dffs[2]~q ;
wire \dffs[1]~q ;


dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[7]~q ),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(\dffs[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[6]~q ),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(\dffs[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[5]~q ),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(\dffs[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[4]~q ),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(\dffs[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[3]~q ),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(\dffs[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2]~q ),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(\dffs[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[1]~q ),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_8 (
	dffs_0,
	dffs_1,
	enable,
	dffs_7,
	dffs_6,
	dffs_5,
	dffs_4,
	dffs_2,
	dffs_3,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
output 	dffs_1;
input 	enable;
output 	dffs_7;
output 	dffs_6;
output 	dffs_5;
output 	dffs_4;
output 	dffs_2;
output 	dffs_3;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffs[0] (
	.clk(clock),
	.d(dffs_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(dffs_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_1),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_7),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(dffs_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_6),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(dffs_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_5),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(dffs_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_4),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(dffs_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_2),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(dffs_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_3),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_9 (
	dffs_0,
	dffs_1,
	enable,
	dffs_2,
	dffs_3,
	dffs_4,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
output 	dffs_1;
input 	enable;
output 	dffs_2;
output 	dffs_3;
output 	dffs_4;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffs[0] (
	.clk(clock),
	.d(dffs_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(dffs_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_1),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(dffs_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_2),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(dffs_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_3),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_4),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_10 (
	dffs_0,
	reset,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
input 	reset;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs[31]~q ;
wire \dffs[30]~q ;
wire \dffs[29]~q ;
wire \dffs[28]~q ;
wire \dffs[27]~q ;
wire \dffs[26]~q ;
wire \dffs[25]~q ;
wire \dffs[24]~q ;
wire \dffs[23]~q ;
wire \dffs[22]~q ;
wire \dffs[21]~q ;
wire \dffs[20]~q ;
wire \dffs[19]~q ;
wire \dffs[18]~q ;
wire \dffs[17]~q ;
wire \dffs[16]~q ;
wire \dffs[15]~q ;
wire \dffs[14]~q ;
wire \dffs[13]~q ;
wire \dffs[12]~q ;
wire \dffs[11]~q ;
wire \dffs[10]~q ;
wire \dffs[9]~q ;
wire \dffs[8]~q ;
wire \dffs[7]~q ;
wire \dffs[6]~q ;
wire \dffs[5]~q ;
wire \dffs[4]~q ;
wire \dffs[3]~q ;
wire \dffs[2]~q ;
wire \dffs[1]~q ;


dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[31] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[31]~q ),
	.prn(vcc));
defparam \dffs[31] .is_wysiwyg = "true";
defparam \dffs[31] .power_up = "low";

dffeas \dffs[30] (
	.clk(clock),
	.d(\dffs[31]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[30]~q ),
	.prn(vcc));
defparam \dffs[30] .is_wysiwyg = "true";
defparam \dffs[30] .power_up = "low";

dffeas \dffs[29] (
	.clk(clock),
	.d(\dffs[30]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[29]~q ),
	.prn(vcc));
defparam \dffs[29] .is_wysiwyg = "true";
defparam \dffs[29] .power_up = "low";

dffeas \dffs[28] (
	.clk(clock),
	.d(\dffs[29]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[28]~q ),
	.prn(vcc));
defparam \dffs[28] .is_wysiwyg = "true";
defparam \dffs[28] .power_up = "low";

dffeas \dffs[27] (
	.clk(clock),
	.d(\dffs[28]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[27]~q ),
	.prn(vcc));
defparam \dffs[27] .is_wysiwyg = "true";
defparam \dffs[27] .power_up = "low";

dffeas \dffs[26] (
	.clk(clock),
	.d(\dffs[27]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[26]~q ),
	.prn(vcc));
defparam \dffs[26] .is_wysiwyg = "true";
defparam \dffs[26] .power_up = "low";

dffeas \dffs[25] (
	.clk(clock),
	.d(\dffs[26]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[25]~q ),
	.prn(vcc));
defparam \dffs[25] .is_wysiwyg = "true";
defparam \dffs[25] .power_up = "low";

dffeas \dffs[24] (
	.clk(clock),
	.d(\dffs[25]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[24]~q ),
	.prn(vcc));
defparam \dffs[24] .is_wysiwyg = "true";
defparam \dffs[24] .power_up = "low";

dffeas \dffs[23] (
	.clk(clock),
	.d(\dffs[24]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[23]~q ),
	.prn(vcc));
defparam \dffs[23] .is_wysiwyg = "true";
defparam \dffs[23] .power_up = "low";

dffeas \dffs[22] (
	.clk(clock),
	.d(\dffs[23]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[22]~q ),
	.prn(vcc));
defparam \dffs[22] .is_wysiwyg = "true";
defparam \dffs[22] .power_up = "low";

dffeas \dffs[21] (
	.clk(clock),
	.d(\dffs[22]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[21]~q ),
	.prn(vcc));
defparam \dffs[21] .is_wysiwyg = "true";
defparam \dffs[21] .power_up = "low";

dffeas \dffs[20] (
	.clk(clock),
	.d(\dffs[21]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[20]~q ),
	.prn(vcc));
defparam \dffs[20] .is_wysiwyg = "true";
defparam \dffs[20] .power_up = "low";

dffeas \dffs[19] (
	.clk(clock),
	.d(\dffs[20]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[19]~q ),
	.prn(vcc));
defparam \dffs[19] .is_wysiwyg = "true";
defparam \dffs[19] .power_up = "low";

dffeas \dffs[18] (
	.clk(clock),
	.d(\dffs[19]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[18]~q ),
	.prn(vcc));
defparam \dffs[18] .is_wysiwyg = "true";
defparam \dffs[18] .power_up = "low";

dffeas \dffs[17] (
	.clk(clock),
	.d(\dffs[18]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[17]~q ),
	.prn(vcc));
defparam \dffs[17] .is_wysiwyg = "true";
defparam \dffs[17] .power_up = "low";

dffeas \dffs[16] (
	.clk(clock),
	.d(\dffs[17]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[16]~q ),
	.prn(vcc));
defparam \dffs[16] .is_wysiwyg = "true";
defparam \dffs[16] .power_up = "low";

dffeas \dffs[15] (
	.clk(clock),
	.d(\dffs[16]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[15]~q ),
	.prn(vcc));
defparam \dffs[15] .is_wysiwyg = "true";
defparam \dffs[15] .power_up = "low";

dffeas \dffs[14] (
	.clk(clock),
	.d(\dffs[15]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[14]~q ),
	.prn(vcc));
defparam \dffs[14] .is_wysiwyg = "true";
defparam \dffs[14] .power_up = "low";

dffeas \dffs[13] (
	.clk(clock),
	.d(\dffs[14]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[13]~q ),
	.prn(vcc));
defparam \dffs[13] .is_wysiwyg = "true";
defparam \dffs[13] .power_up = "low";

dffeas \dffs[12] (
	.clk(clock),
	.d(\dffs[13]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[12]~q ),
	.prn(vcc));
defparam \dffs[12] .is_wysiwyg = "true";
defparam \dffs[12] .power_up = "low";

dffeas \dffs[11] (
	.clk(clock),
	.d(\dffs[12]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[11]~q ),
	.prn(vcc));
defparam \dffs[11] .is_wysiwyg = "true";
defparam \dffs[11] .power_up = "low";

dffeas \dffs[10] (
	.clk(clock),
	.d(\dffs[11]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[10]~q ),
	.prn(vcc));
defparam \dffs[10] .is_wysiwyg = "true";
defparam \dffs[10] .power_up = "low";

dffeas \dffs[9] (
	.clk(clock),
	.d(\dffs[10]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[9]~q ),
	.prn(vcc));
defparam \dffs[9] .is_wysiwyg = "true";
defparam \dffs[9] .power_up = "low";

dffeas \dffs[8] (
	.clk(clock),
	.d(\dffs[9]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[8]~q ),
	.prn(vcc));
defparam \dffs[8] .is_wysiwyg = "true";
defparam \dffs[8] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(\dffs[8]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[7]~q ),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(\dffs[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[6]~q ),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(\dffs[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[5]~q ),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(\dffs[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[4]~q ),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(\dffs[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[3]~q ),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(\dffs[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2]~q ),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(\dffs[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[1]~q ),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_11 (
	dffs_0,
	reset,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
input 	reset;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs[39]~q ;
wire \dffs[38]~q ;
wire \dffs[37]~q ;
wire \dffs[36]~q ;
wire \dffs[35]~q ;
wire \dffs[34]~q ;
wire \dffs[33]~q ;
wire \dffs[32]~q ;
wire \dffs[31]~q ;
wire \dffs[30]~q ;
wire \dffs[29]~q ;
wire \dffs[28]~q ;
wire \dffs[27]~q ;
wire \dffs[26]~q ;
wire \dffs[25]~q ;
wire \dffs[24]~q ;
wire \dffs[23]~q ;
wire \dffs[22]~q ;
wire \dffs[21]~q ;
wire \dffs[20]~q ;
wire \dffs[19]~q ;
wire \dffs[18]~q ;
wire \dffs[17]~q ;
wire \dffs[16]~q ;
wire \dffs[15]~q ;
wire \dffs[14]~q ;
wire \dffs[13]~q ;
wire \dffs[12]~q ;
wire \dffs[11]~q ;
wire \dffs[10]~q ;
wire \dffs[9]~q ;
wire \dffs[8]~q ;
wire \dffs[7]~q ;
wire \dffs[6]~q ;
wire \dffs[5]~q ;
wire \dffs[4]~q ;
wire \dffs[3]~q ;
wire \dffs[2]~q ;
wire \dffs[1]~q ;


dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[39] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[39]~q ),
	.prn(vcc));
defparam \dffs[39] .is_wysiwyg = "true";
defparam \dffs[39] .power_up = "low";

dffeas \dffs[38] (
	.clk(clock),
	.d(\dffs[39]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[38]~q ),
	.prn(vcc));
defparam \dffs[38] .is_wysiwyg = "true";
defparam \dffs[38] .power_up = "low";

dffeas \dffs[37] (
	.clk(clock),
	.d(\dffs[38]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[37]~q ),
	.prn(vcc));
defparam \dffs[37] .is_wysiwyg = "true";
defparam \dffs[37] .power_up = "low";

dffeas \dffs[36] (
	.clk(clock),
	.d(\dffs[37]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[36]~q ),
	.prn(vcc));
defparam \dffs[36] .is_wysiwyg = "true";
defparam \dffs[36] .power_up = "low";

dffeas \dffs[35] (
	.clk(clock),
	.d(\dffs[36]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[35]~q ),
	.prn(vcc));
defparam \dffs[35] .is_wysiwyg = "true";
defparam \dffs[35] .power_up = "low";

dffeas \dffs[34] (
	.clk(clock),
	.d(\dffs[35]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[34]~q ),
	.prn(vcc));
defparam \dffs[34] .is_wysiwyg = "true";
defparam \dffs[34] .power_up = "low";

dffeas \dffs[33] (
	.clk(clock),
	.d(\dffs[34]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[33]~q ),
	.prn(vcc));
defparam \dffs[33] .is_wysiwyg = "true";
defparam \dffs[33] .power_up = "low";

dffeas \dffs[32] (
	.clk(clock),
	.d(\dffs[33]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[32]~q ),
	.prn(vcc));
defparam \dffs[32] .is_wysiwyg = "true";
defparam \dffs[32] .power_up = "low";

dffeas \dffs[31] (
	.clk(clock),
	.d(\dffs[32]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[31]~q ),
	.prn(vcc));
defparam \dffs[31] .is_wysiwyg = "true";
defparam \dffs[31] .power_up = "low";

dffeas \dffs[30] (
	.clk(clock),
	.d(\dffs[31]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[30]~q ),
	.prn(vcc));
defparam \dffs[30] .is_wysiwyg = "true";
defparam \dffs[30] .power_up = "low";

dffeas \dffs[29] (
	.clk(clock),
	.d(\dffs[30]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[29]~q ),
	.prn(vcc));
defparam \dffs[29] .is_wysiwyg = "true";
defparam \dffs[29] .power_up = "low";

dffeas \dffs[28] (
	.clk(clock),
	.d(\dffs[29]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[28]~q ),
	.prn(vcc));
defparam \dffs[28] .is_wysiwyg = "true";
defparam \dffs[28] .power_up = "low";

dffeas \dffs[27] (
	.clk(clock),
	.d(\dffs[28]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[27]~q ),
	.prn(vcc));
defparam \dffs[27] .is_wysiwyg = "true";
defparam \dffs[27] .power_up = "low";

dffeas \dffs[26] (
	.clk(clock),
	.d(\dffs[27]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[26]~q ),
	.prn(vcc));
defparam \dffs[26] .is_wysiwyg = "true";
defparam \dffs[26] .power_up = "low";

dffeas \dffs[25] (
	.clk(clock),
	.d(\dffs[26]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[25]~q ),
	.prn(vcc));
defparam \dffs[25] .is_wysiwyg = "true";
defparam \dffs[25] .power_up = "low";

dffeas \dffs[24] (
	.clk(clock),
	.d(\dffs[25]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[24]~q ),
	.prn(vcc));
defparam \dffs[24] .is_wysiwyg = "true";
defparam \dffs[24] .power_up = "low";

dffeas \dffs[23] (
	.clk(clock),
	.d(\dffs[24]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[23]~q ),
	.prn(vcc));
defparam \dffs[23] .is_wysiwyg = "true";
defparam \dffs[23] .power_up = "low";

dffeas \dffs[22] (
	.clk(clock),
	.d(\dffs[23]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[22]~q ),
	.prn(vcc));
defparam \dffs[22] .is_wysiwyg = "true";
defparam \dffs[22] .power_up = "low";

dffeas \dffs[21] (
	.clk(clock),
	.d(\dffs[22]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[21]~q ),
	.prn(vcc));
defparam \dffs[21] .is_wysiwyg = "true";
defparam \dffs[21] .power_up = "low";

dffeas \dffs[20] (
	.clk(clock),
	.d(\dffs[21]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[20]~q ),
	.prn(vcc));
defparam \dffs[20] .is_wysiwyg = "true";
defparam \dffs[20] .power_up = "low";

dffeas \dffs[19] (
	.clk(clock),
	.d(\dffs[20]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[19]~q ),
	.prn(vcc));
defparam \dffs[19] .is_wysiwyg = "true";
defparam \dffs[19] .power_up = "low";

dffeas \dffs[18] (
	.clk(clock),
	.d(\dffs[19]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[18]~q ),
	.prn(vcc));
defparam \dffs[18] .is_wysiwyg = "true";
defparam \dffs[18] .power_up = "low";

dffeas \dffs[17] (
	.clk(clock),
	.d(\dffs[18]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[17]~q ),
	.prn(vcc));
defparam \dffs[17] .is_wysiwyg = "true";
defparam \dffs[17] .power_up = "low";

dffeas \dffs[16] (
	.clk(clock),
	.d(\dffs[17]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[16]~q ),
	.prn(vcc));
defparam \dffs[16] .is_wysiwyg = "true";
defparam \dffs[16] .power_up = "low";

dffeas \dffs[15] (
	.clk(clock),
	.d(\dffs[16]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[15]~q ),
	.prn(vcc));
defparam \dffs[15] .is_wysiwyg = "true";
defparam \dffs[15] .power_up = "low";

dffeas \dffs[14] (
	.clk(clock),
	.d(\dffs[15]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[14]~q ),
	.prn(vcc));
defparam \dffs[14] .is_wysiwyg = "true";
defparam \dffs[14] .power_up = "low";

dffeas \dffs[13] (
	.clk(clock),
	.d(\dffs[14]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[13]~q ),
	.prn(vcc));
defparam \dffs[13] .is_wysiwyg = "true";
defparam \dffs[13] .power_up = "low";

dffeas \dffs[12] (
	.clk(clock),
	.d(\dffs[13]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[12]~q ),
	.prn(vcc));
defparam \dffs[12] .is_wysiwyg = "true";
defparam \dffs[12] .power_up = "low";

dffeas \dffs[11] (
	.clk(clock),
	.d(\dffs[12]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[11]~q ),
	.prn(vcc));
defparam \dffs[11] .is_wysiwyg = "true";
defparam \dffs[11] .power_up = "low";

dffeas \dffs[10] (
	.clk(clock),
	.d(\dffs[11]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[10]~q ),
	.prn(vcc));
defparam \dffs[10] .is_wysiwyg = "true";
defparam \dffs[10] .power_up = "low";

dffeas \dffs[9] (
	.clk(clock),
	.d(\dffs[10]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[9]~q ),
	.prn(vcc));
defparam \dffs[9] .is_wysiwyg = "true";
defparam \dffs[9] .power_up = "low";

dffeas \dffs[8] (
	.clk(clock),
	.d(\dffs[9]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[8]~q ),
	.prn(vcc));
defparam \dffs[8] .is_wysiwyg = "true";
defparam \dffs[8] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(\dffs[8]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[7]~q ),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(\dffs[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[6]~q ),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(\dffs[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[5]~q ),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(\dffs[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[4]~q ),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(\dffs[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[3]~q ),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(\dffs[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2]~q ),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(\dffs[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[1]~q ),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

endmodule

module SerialFlashLoader_lpm_shiftreg_12 (
	dffs_0,
	reset,
	enable,
	clock,
	altera_internal_jtag)/* synthesis synthesis_greybox=1 */;
output 	dffs_0;
input 	reset;
input 	enable;
input 	clock;
input 	altera_internal_jtag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffs[15]~q ;
wire \dffs[14]~q ;
wire \dffs[13]~q ;
wire \dffs[12]~q ;
wire \dffs[11]~q ;
wire \dffs[10]~q ;
wire \dffs[9]~q ;
wire \dffs[8]~q ;
wire \dffs[7]~q ;
wire \dffs[6]~q ;
wire \dffs[5]~q ;
wire \dffs[4]~q ;
wire \dffs[3]~q ;
wire \dffs[2]~q ;
wire \dffs[1]~q ;


dffeas \dffs[0] (
	.clk(clock),
	.d(\dffs[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(dffs_0),
	.prn(vcc));
defparam \dffs[0] .is_wysiwyg = "true";
defparam \dffs[0] .power_up = "low";

dffeas \dffs[15] (
	.clk(clock),
	.d(altera_internal_jtag),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[15]~q ),
	.prn(vcc));
defparam \dffs[15] .is_wysiwyg = "true";
defparam \dffs[15] .power_up = "low";

dffeas \dffs[14] (
	.clk(clock),
	.d(\dffs[15]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[14]~q ),
	.prn(vcc));
defparam \dffs[14] .is_wysiwyg = "true";
defparam \dffs[14] .power_up = "low";

dffeas \dffs[13] (
	.clk(clock),
	.d(\dffs[14]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[13]~q ),
	.prn(vcc));
defparam \dffs[13] .is_wysiwyg = "true";
defparam \dffs[13] .power_up = "low";

dffeas \dffs[12] (
	.clk(clock),
	.d(\dffs[13]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[12]~q ),
	.prn(vcc));
defparam \dffs[12] .is_wysiwyg = "true";
defparam \dffs[12] .power_up = "low";

dffeas \dffs[11] (
	.clk(clock),
	.d(\dffs[12]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[11]~q ),
	.prn(vcc));
defparam \dffs[11] .is_wysiwyg = "true";
defparam \dffs[11] .power_up = "low";

dffeas \dffs[10] (
	.clk(clock),
	.d(\dffs[11]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[10]~q ),
	.prn(vcc));
defparam \dffs[10] .is_wysiwyg = "true";
defparam \dffs[10] .power_up = "low";

dffeas \dffs[9] (
	.clk(clock),
	.d(\dffs[10]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[9]~q ),
	.prn(vcc));
defparam \dffs[9] .is_wysiwyg = "true";
defparam \dffs[9] .power_up = "low";

dffeas \dffs[8] (
	.clk(clock),
	.d(\dffs[9]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[8]~q ),
	.prn(vcc));
defparam \dffs[8] .is_wysiwyg = "true";
defparam \dffs[8] .power_up = "low";

dffeas \dffs[7] (
	.clk(clock),
	.d(\dffs[8]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[7]~q ),
	.prn(vcc));
defparam \dffs[7] .is_wysiwyg = "true";
defparam \dffs[7] .power_up = "low";

dffeas \dffs[6] (
	.clk(clock),
	.d(\dffs[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[6]~q ),
	.prn(vcc));
defparam \dffs[6] .is_wysiwyg = "true";
defparam \dffs[6] .power_up = "low";

dffeas \dffs[5] (
	.clk(clock),
	.d(\dffs[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[5]~q ),
	.prn(vcc));
defparam \dffs[5] .is_wysiwyg = "true";
defparam \dffs[5] .power_up = "low";

dffeas \dffs[4] (
	.clk(clock),
	.d(\dffs[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[4]~q ),
	.prn(vcc));
defparam \dffs[4] .is_wysiwyg = "true";
defparam \dffs[4] .power_up = "low";

dffeas \dffs[3] (
	.clk(clock),
	.d(\dffs[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[3]~q ),
	.prn(vcc));
defparam \dffs[3] .is_wysiwyg = "true";
defparam \dffs[3] .power_up = "low";

dffeas \dffs[2] (
	.clk(clock),
	.d(\dffs[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[2]~q ),
	.prn(vcc));
defparam \dffs[2] .is_wysiwyg = "true";
defparam \dffs[2] .power_up = "low";

dffeas \dffs[1] (
	.clk(clock),
	.d(\dffs[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\dffs[1]~q ),
	.prn(vcc));
defparam \dffs[1] .is_wysiwyg = "true";
defparam \dffs[1] .power_up = "low";

endmodule
