// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HUra+O15AO2BgnjiXKJrhcRf32KSD7R5oE+GaciKGXtkDxt39KSpgG5mTtA8QhpU
OdvV3iwxconqO4T/ZXig7ITLBnf8OjHKgg/Cm7vAh6MsSxJuU9cWrcZqfXLwRPr3
gW3OiqJwoi6UPLOVi/dWbQrGzHxz6dDGt332ZijsIMM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 49312)
GICxakIGY+YHIrZ6B4n4IMzLWwuELYBJbeMqILPw6luco8Rxv/gTHJPhI3ywexlw
9BpU5uWouoQIJxmU5/ivklqjM/O0JfrMag4m4CiuJCddOVAf4IjV+T5U51YkrPcs
IBITwMnEGUbA5fVpqWfoxBzilUjregCksbEYFN6I1vtV5BwdlM7DOSUKdhPIVe/l
HSbuyUAJ6Lfzx9MbxyYifLNgOxqYQ705otwy29RlPHAUnPgHACOf7Ggt+8/WBUg4
MzLc/zy4ZgAogcMY9I4dhJQWv50x/iGaykssYoIYXbP/QDBPvpf722CoGMU4U0cc
i8A3eLSZhqYQT1JXn+4NdEO8Ks5Jfj++pt4rgQCmEcgNl55q9tAPsiaF3T1eCI9r
imWKppXAHkhFFhXyL3GAOFSPJnoigTnMLUiRAbOOyVkXjHHYSGqPr68EPh84q1X+
OfF9qG/TBiaag+2st8KA1IIcWBz72ucizYpNGtVSrVm6yHy3MGAT7f16+ytKD3bE
76GnYbC1h3xu0xrtHKHyJR1mr3gX6OstOH1WxFZ2kKTAwDZYWvke9QwfZ1XTPutu
MwtykorMyoHoB3HkxX5uIfJAhw+gexQEAd/wMkCLyG7FCHWdh+7HG/voBU6mkRcH
Eju+Tb4rCk9P5yTRdKItyfq16ztVeFjC58DgZ4GWUGR/FrnbsNcYO9ZAqZQsUUY9
lUVHR1d6G5gsF6qNcf8ZrSovbYsIUUDJOZfCxMm0wONAsE4Gy8KG6zzIPZPtnFZX
G2L7aW5zC7DRp0ZT7rP4DJ57ogYv6y4hs9360xM4VGc5ZglKwNjuhUxEykzBMopk
UD63Hm3hnpm6wNH8wuIBVzE+OHpAGllEoAcTT3+K+bmzF8OS9KUgq3V4ajZbih5F
XJfNrOy/t95vNQce+Vf4y/Wf/fkqhvJuVUBSp57dlpcCKT8EOq66pp3roch3vxo9
E3nGtJ/4DSFh9ZTYiGNEru4wAbGpV1dkyPcOmtsqeQ5q/sR+3D1QsCaWhEQSot5g
VWtnEPCDbo1qpYw+ADaopCK6udyUjcBhim/2nXwcw5PB2/eapIxXh4HgjoVSJBuw
RbizvEkndufI7L/qtmI6OVe7q8IIhTe8tR4Vbn/KG0u5aFo32H8qGtiiqrINyxZC
+SbUM2l9yHr6jdfLau/NNg6ux9e8b3/gxKMVQiw5sY9DiJv5Vep30JjogpFl11ul
CEmycrqDQK49OJfmVZ/9clvnqxNOfH9stJe76YnK4qba1OmczEDQLYWQgygYW1GY
B1jvBZTRn4Rl/4jOMXwO63oNq+xFyGTRPTSFlye4wdV/B7aNbkPxHjGFADfRWele
Qu8YQ3pkeqXTUgCk6yb4/zXCynUGuw0WRx0tGko0Oo4DAayTdksKZYC/GIt4JIa8
KPwBiFGzFHz7Ek5cUbsfithUa+MQyZKtWqlZu+133PYrrNvZl0JfHTbxwlNC2JMQ
D+XUo8FEXSbZsFLyeeLo7dtpxc5xkxcxQfz4vIHfgSUUS9S1D5XMAwWMAs74GhbV
Z7YC6HjW6+iIQ1ogkXSEtynmNATqeUX2qtAmjh33exP8J9xY2vc6OrI+n0HZ5m6Z
/VLUtCyCPLl1YqK1bLLk7RZOlmKcRq1kJYlSf/N0PUBCV7633xeitdfGgf9N6QFj
a8hXBYsTny5Glc8gs4gVn1ykpf2X/DvwqT+sFOjpJ05KUbZ6satoSHy3hel0wGV3
LmkSApAhqhtN+nyN2wr0bskoVV1d6/urs1Sky1z7En3pG5Zc+sB/9wa68pbVQmne
Z3x1EV5L0RGwlUSrUoqPBb/bT+yaPqVgM/A9boLvQ1mGdH9bltSoLUIC+YsHTSLe
bQENOvKFlD0Dryx+NOgs3DQuIaTYVuLuiNiUYcwS4U4ROzRMefinrpt9imbJcJMt
BCjrJtQenTZxDRaTt6BmvqMVRnXZOmh/SnWYTcwWZFIbkqD/yXpJzInPKy7oY7nE
FuUNE8XmNrKQis9+PjwllccQXjMi6fj1Uqll3oRwpHdwNxOB1Kvpravia+D0puuK
d4I9SJTXbkKP2WlKCnMWxW+/5xgOGOQNhO8R/e8yK4x2jX7kHL5g6UtZKHV3zCF+
KAiZAAQahyZZPNIt+6uc+3DqgX33l/GOQ6nUDHyZZJahLyaiMq2jW/iMSO8taE1o
3bL0nsMjbe1Yv9GgehQYOb5vn+hNkC9oio7171JEp1gb0Q3BKNmvnWJd8l6o2DA2
/oKNv0kWfHlqLWBViroVy5kPaCPF+FvlH260xUnmfKMGeCAxJHflKPrN7XDgxQ5K
8nIJwgxN6KOyd9ShN6J+Pv8gHHP69eQQKwUa99bAIUds0p7N1zb9vqLGliZCj6dM
WfIFfMMYQ8ulZaMWMYIU5zJDEQ7zS1iJvAIo5ru49rq358gstlb0b8eshJaEQd1d
x67sRiC32UxRMR3YGCT7wIySUe0rfOS2vyjSg0f7ZtYgpCux5yeAgFpTk5HxDLzN
oyV4mTAw2SZOblHXOSZcqT5SYO2WUF4MNNTiHVz5S3Q6+sEJi9ZqBfoFgts/9wBj
l0f58QyFgKF9sBD3f54yCz78VgRcUno/mr+M/Z0G3ya4FMmtIp3cojJNq1OrACnL
s9YnvuJf35VhATbQ5squj82jtZVpVrR6Ng4+5UnW0uMbmuMyw8RKtNCbowIRTM9C
qRrKzR6ER4hlU0sPRcIhbXjXgM+xmSecs2Mqk1wrFXdK5ZVFgBrRCUgq6UYv3d8H
aO3kVatOF441tRL6G9IKl64H7qkyE4gOKqD7JOIIXY1WiXc4wpUUoKg1/0Rwp3JT
KELM3bPeEt3r/WqneBQcRWYa8Oqgs8jUgCwKFXSZ7seNxVlBwGyhRv/F1Neiny/N
NMyEkmN+6dPUJiWseNxpzd+x9EvxbJmqQWBogOo2fUDmftMBkb4clSLvjXM/iRVx
Alf5aEWTtFNosbay4XWVMXP5MjvQwuSHiCLqtwfV4SHV2YqP+o2BxMA9Dz4//Kvc
KDYILraCWLomZM0BUMAlxwukbsb49CwJO7y8YIRoY4gkySKAUYO/7aLFy1CYpK6B
0D/PE7z7zgW4zRHl7TT8zOLxPKVCQmLVPYGLzpj/wI2mZnp5NKEQ9SHUqLd+VN5h
sJnEJtxvu1qNb1Q3+VywYNuUFy/vA4jAYZPVpxXiuGaW4QrDVN7YaO5iy4JU1PoK
cNnq2D/bjODwUB3v77sSqZexnfm/YoM+2QtlVBMwhaH53smp3Ju1p6l7e9XCzmUd
/S5N/QCdPYHMtsXPjH+CUK6ztL9Ez6VE2tboY4saVoto5LQpYk6QR3FbZcfkUGP1
ndnEiVUe+2nlDBM1rff1AroK8FASyIelfVZrzQ2Q+vOlfg4zHOPmGBUOMramAnYD
brGklYvKr+kDxMDdUmcdRoWtq+N4K3KO/KJNmHXmWpfRA9W6D8W2OqhvKdI39CfG
DYghp/xXIgtXm6lLSxfDVWsxZGfX1j1PxQqE6ywsDb3JWG7YN0sy/Q9AHrMHMC9m
RroC9JNruApOTnFMv18m8vahxpp0U5pHAz84BjjYETivsiEIUeyd+TvNroLjrDTU
Y2c2EaUxkSROSTCHOODZCeHxSRrrmRX01Glo9A0EhUTbP4ozQq3zyh/yJUt+FmJS
7l0NmYyT6noHlqwQF4961FipJDrGNzut/tC9cgWbOU0B+DBO5YJubWTXK5e9jJ43
+3lfypk5WI6ln0mKA+OlpFS/4q5BhlakLhM3QXpgNaqM7QGhg0/6yR9uzm0c9yWF
SifxBlLMPeFPDUPWw2Reoq65AwMoezd7EWB4qpNqdXIqEtQ7cXD1U1KgqpSdeyFq
eG5oaYrSXSF47lroXnP3S3XIqchqh99TtobQY9otGX/LoYUxgj86mMoiW3JJ6u0/
nQ7Ij4FEDglC+mLhN6frx7Huhc6vWIji6T7x7Pldetyvwby9lEjfnRdveF2mrSLN
N4kp49At9kFwKdBkxV9jEbWwiCW9lCLeh5dO/pR1NQsPiW+CN9f3j3DruraWF1Pl
hpv2XlXduagf7MbNSXtSKRyIIFVPVTNwZH0stbugh4LGnTrmyvQl88G3w09a2bIf
gdviGAIPIFYoJaczb9h/KNUXWsFrp74vvTNuDyc0I/+lN6avjUccbks0JP3vVEPu
grQDXJwsqQy+sCw5iqUMCARBLxLMNAJib3Y7NYxGmE2uVhYuvgrJttbaqHAw5XDY
DJJMLTuW4WzI86+rRmVE+8YCHNltlDpt5HiJJKpY86zljPZNcuXEp4bf4+26DOm8
9zMfJ9pbuhnx7sTIJ9m4Q5Fv/TviXpWozZCFKrEObEbwfA3k46Ts/nq8MTIi68vw
HJJwsdHQViULZ9YW3PbTuUwYZ90N2BTnwJK6E3AUyGVCTxd9MQAmmZY1bG4UHLXP
orNtl52Fgvh+r3Ek87D0m2XoPAWY/HZCmcXpvylh23dN5gKKS3rKGkBRuhqLsTLB
4lMvT03HHy3xF3JJir15ZTrs42cHK3FaHifIF3LcN7vwfsG1r9yM3Wa2HsbUPD4N
GLTQz41Ls5h1ol5EYd8+l/ljFCqoaWL1uERx31VaFywM4bCdKzF/XoGBaCo4uzAO
tb7J/6GQJh8UvtoxtUZn/8lts6KfoG1ypT02NAuuwjYXI6kXEwYIYOijr3BcHmj7
9TJFWsJzN0SHhmZxhhYvfC3h8ieOY6TNY0R4/wKaCvyrDaRUSDSfWPj3S6VOyd4O
MlZLGf0cK+TT45kGnIV0/euKj1coCYVmQr0UCpLRKaSCZF8UyHIpqPDUSH/L0/TB
IgJSLV++s1SFq9gWzCGJULL/ZV+m7HJAQhPj0IZSWLKi5z/yuHaQHplW9hfl3W+M
9UAJ9JDnsdwNBbWF+QnB0sa6kyUOUDqEzgtMLSQ0pcNthnN3CgiWqZLALyvmJHiM
4McwHAOWdWOmqsbuPdXV+YYXQ7h37f2XJvirvo524zXI2+Tk6v4aANbbgohSMxaO
BjEyvYyRLNHzEsIvw/8xHVa636KHniApyi+salCfgWkY5YyTlDzok/ABSTGMzjPy
Ovc3mN3gG4E+bkoKeSgxxIDz+0+P0/h/5voPdGyiJb6v09MnxhC21wFjExWEZoG+
AVNkPGaYaLoBKqpoQmidvtK7s9WZFsQY2nLvzJRZP1j0bPcmuIb5dQWEEU2LlxUR
NZLGBSDU4OhRxUbg86n+Z+TLc+HVLcYcxcMF8Gj5xTMmDFA1DRi4XBPY6jbtajcs
DOez6ebtS/t81IZYmCYwcNwYPj/OH7PoXGE9BPdunl+PAOAwH6kbcryn4BkxFbLo
qt8Q9Q+EhTjSUe6DzthanthdMpC5w1usi9hL7A54qTkEEyUqRB2oulV/XGTaca1z
voXdJr+Gsvz6F8XriOtUGLiySv5OeBEqdHuRtkjQsI3bzRXxx8voyotkjKqlGkr4
gMzlXj2bL8U1WJm+KDTMlFVt8wMVAurmDF4+YJmV0BGEMCk9nQ96p3det2zXRgdq
Cy/L6gU76UI/lQ4cCt9j42v46fl4zzTQgoqMLe4DN8FAOr3E6i8ws1AFwyGh4ihr
gMQWVakT7P9QTS3HPRwFC3WBCU3nVBpTBK5DghKhCqka8KKSWg05FCgLFo7gSYgZ
FQKJKInX1JUF13U43R+RhTqtUENeU7427twdAwvBix/9WwNjip6d1LqBh2jgcmZx
r2tTNDCwmXmSFQDVNGcFnCfTVS6E+RnvZk7A1xk4/xKDHDcGu351puwrILhHcgSU
2Il8RwplBsm8h2iWuysae14OFacgZvf9CP/C7aMbGU3Mpdh0wxaKbidq3pbTXPDi
bHMt1TNy0XNORwtCrK8K9PPWiMY+D3UiNZsdKwxcKJeCbHPedRTnhOIm3htdMBql
iSsiA96OYldXqc2SD6Qgdcyv3SuZfTjnQ/mtqvGusfe9LkWD/wqRA2nJ4ee8NnW9
uEqR9iSg6xvLjvHZXcn+tdeN+bfRnarZ48VcBAyTT207ELaycoWBFTGpcraA69z4
mX/9AI3h+lbuFs9sPorQDUI7ARXNP8cXXRusXZiEgEVxccO9zMN7Q/gLl1v/w5HB
rBJRjBdr5jHw0+ycoUG8V84vYERBmVf+mKXDyhvviv1gr+E4jJe1gI6wuHNykomH
6fLIJpoiHtwEDCCkBiSLanFPK/ZHC6EVuyEub81Ux/9R4UUBn8OlEdXtiNlL+Pkg
oWGRH9myYN9NFKEDFOs/PtYsQvHRsOrWycNbf9exG5HdLSsR5qtlCdyE4WnQfZ2x
FephFnl9l5CDWGLc0ABSCCVRkB5mYx0Ur86xgqGBOVegxr4mdHD8vSBJ42iQBHDM
6aGqS/8OI/YM79Ne/g8Xwj2fEZgpLcLU5mKZv/KoRpgDvjxjAY0XmAwsoqeMILlC
LekHWkzflR2CCX6sb+U/fclspePzmQFze+zf1rgjTkSCXKzox7LH6o/3o78Oj1VV
IP7XrByEOmE/yJM8YoYqVfsBjdnS8ohjXW4Wvc4r0cd0WM7QI6CtMTxwAJO8z3ao
x8S0Qv2bCWUpw80Bvy9tlnK8GHL1ltvhyhH0ZkPZliivSu6k72Grf+NrklFCQXCK
ouio5o1dd/Q8M67viHai6ud4OdxLhhKQEt4+x1TUrCVslxOcoBY+R8GefLcucgfK
WoXpzA6uKc4FXLkFZmrm+eCsBS9dL9BZgjxvw/sph1yHHZXW4TF0p78PA7M++s95
tvp7McU6m4CIeWK1LeHUkeivEmUN8WzyHf9kifCLymvcouMrzfMY6bSHrc6vPr8a
7GIAQT/KMViwsaOjtxPBgctoHsnRINKeYOlTMhf8wT8tASTCRoHJblz8vCY0WqGI
A/vZfRAQMXhKd4Eq7FKob5IQWpcBQewV2wFBm6F+AtYZzTrPBNp/KIM0ZGluTD3x
1f9gMXSoNVGFjEIe68fjCAD2wlk2Ne/omezCIteCCpqXT6j2GbIZ92ilnOHjjOk+
D6j3phLW/3WWeSEARvJznpjSch12GgEqpKkmKNLKIyh7qGTNHoTtGAnZxrzDqj82
V5qYEmuXZXgdxF4Zeit1dY1veu32x4SyFHM9Bq7InBdhPsIl9112vfkjgEEhKBnB
jQpm+AKmB9zz4NQQdn2HlanE9pQId7uKr80+CHwGam8IWVO1W6slifZDOtMnEMnc
myk7xveYAs3JhBhNmVn6VzBR2WAxyW5rBUFg6y5jVYeQP2lN5+pw43dFE+LEPHZV
P9liULfM6VcBXId8O9AF1n7gpSuFIZbR07dVQ8PnIsISpMR1UXFWPWXjMMDcFpWq
3d+YzjImwPcrjDe8fYY+6NKmlrwILoz3M7rp0S0VZS1mCDkuS5R5aGQR4rk8PRnk
N9tMO5fKTwcG4TynbI3FpCZTTVOB0IHLCmJtxRq6wijVL+pWqMYR0egG7yURIPMf
mZy08vIto+Sq0qZ94yRmQlbmPHztR70QgOX7R7qc5tNaywRE/4iZaNGvdg1wgyn0
8zlRANmjmrLyOdY4uldgv3xrRk0NSrNGZQbG5Qx2r8IpA8GB8sF+PAS5d/CxVR4+
h2dYMHfh9cLwNvZkVPqqdCdc/1xes08UFqFIlJt4+5fO5aDacMG40PBuKRhHrJ1t
tjNdfyQ0YQ0d0RbyINrSR6unAA9SxccFdtzLCUrZk5bTMXq4e+PDaNiEhkxWjjq0
mXgdtV4LVmArkMT28NltGZ73MImYg5ol8t8v9sN+vlY7+5Z0QcThewtekTlVxgdi
JDaZVS4Z/jsXL9v4WRIf6hxUBK9zf94ApNTKcbA0efZKrtot1h0H9zvJp8fk5oWM
yyweK1Kc1h6iT5ipEl9GZ5U/Pl7+qs4lXOz/uY5Iwtce69xjWQCJzpzLGOUZ3UMZ
0kIRPTxv0I89AA6v1ZgSjsVkScaH9jgroGCAnqHK9X8mkem3NbAQuzzbd48Q896B
L/vTiMW4bFs6AD4SOGSdGfLQcjgJoG5y42ftMf8dmiOPGu5HYfblCT6kWY1X3nBK
YOhJQacT9Oh3HkmjoVZ1qaSY7gDqJYMi1YTuvbdZbrMpJriD9y2YwL9eOMeQ7w0p
KRLHhG6TzP+frN1Fw04miXHVPvV7purI2oLc1aT0xCENTcbcjVPM38jX6CsP0Kq6
dhDphNM/R/ulGrI/yWPtbG6UYIHErCQjTMmsCjqS5O/Gx0SHGlub1VjwxMj/5dQB
ug8h9Mol8cNibVEubRJeX+jqEIgfezplJikxeAVse1n0MeeRLlmIZZPySPXikfxk
dA+E3FnnbMGeIQ56Aw5g6GYK3bamv0r+PNDpQGDBi337C3RH6yWl4f+j+ctcZX7p
6SNn+dH+5md1uUqKQbAsrgj9M8WZHrpAUSzEAnND5W1J+Hltt7ePLDCbgrm93gZw
esCgM+0PmTSgJDrk03ud3WcM6+N1w3+8wdXnMdFqKf32cE5gflPKLPw+vSCwTvzP
3gB7TbaBjv+n/Q+DVJIwKv6hi5plLpMPlAoc5gTwng8SP3j3RXamLbIYwPGg94zI
9QpTavjF5b+sAzN7k8huNM6oydt3ScanQfEAem/1sw0cg6MjTjbg1fx9EmjWmj5P
EpYJ/t9ZRWUTVfRrwbnohdhhjaroOJ2UgR4sNuLrsdbQp3w6BX2EEy6Ks7ZLKk7r
aIl+gpQaKVisTHfwxlcG6shn7fTFQsWL2A7LEixNrCkyPUywi5RdTCViBPhjqa4R
nIVdsqsvtoxzYn0lYxe4cai94SeE5rjVCeNARw4Ut9OH3svUn0VAi3pF/c2bBeLQ
UZDw0gIYIQmXKjieXzCrUJIhH+UNtVEKsjft0+L0OP+ABRNs3jOLXd0KQikmrgPr
QkywYUBqvha8jj4lTQYbo8lWDJPXzVb1UJnlj04Wot5kcuLeqIWTQOZRnRCtaCZD
vAgRy6EZZnN1c0/uUv3G/ky+CHF/n90elym9GZ//yiPszcqXneGGgREV3b1EREjJ
C8SflCyu04+6VeaPysVeJZ3xoAymGGvgUyOin/VHQ71OqeHLyBXhKgB4F/VIvSn3
5DfJx8JvPR9f3qOzu9ZfcgC6dmfi9B52Bp/dUH3yTf+CDkxK7ZV2ShJsAOYrwyJD
uXDihfKWxvl63HvLewX1FAufdIRidTJSJEASYmJDS8pFWYRUjTj6qxTilkAF3MoK
0+Tn1/uLB/cXYM1KiaYQlwTXQLdBJB6d+PfHpPPW4uVfaHhRxPSQokg1qc9i5rx2
8xgtlLVt8Qp/DO4M0YT0kuqjgZPXzmkbBXP8MBFRz3qpfVChkMzqzCTyYcl2fAC8
DRaIJtqDHSwUMf+JcwzupxPxz2iiZjy/Oo8OvWsdyYZShbYC/8SinBrYS9U+yJiG
gEQry7Ou4k3VRJuIfkeU3BEI2Ptv/OZU0nUkN3rqa9iPI2cenJommJx0Tj9JfG1K
xD1LjkcGNkq5IjI1rzgK/MYJcog1DutKQGNyDikVkVdq9osVKxTa+aBhyKRD4Fm+
YafhFNhTBa+rY9NzRxqVz6HGomX0aUDy37ZZf04SXIfIM9qUkLERH722l9fGDQgA
S47SP6jmrjXgBgJ5MOi9t/Saa7wVmMVbeMtVfoJS8w/7uqgwV2ud5AtLsstwQTpJ
FdQE7Gty7EA3hGQRvDnKiI0Owk+6CUMByqObLmUd+9ehrrB5gxgO9KH8VPAcD7RU
XdwuNuy2U9yGVlM6Mo8gOHCo/QUGMPqlHMfDtBNi2DlpaAC6JWp7tW8q/fd2nfcy
5HGtMTY2c08T+pWkyTs0ApdJWznBHxdXfxgvL9IfCld7+bvAojysj+ylC27iwHdz
UwL1SyxK071XwSO0HLvjSG4I9N2SmcLK01heJLj0mjOQM5xEJWy88jaA4i50cg+v
n0Rol8MPRhCCXMg92XLhPIFnW0crX1LAtoShXC9K+TyKum+y93vBn6znxnxT4+Zl
ZSnMsO8ryp1YnClUX+o+z9K0RPT0D3XLbb1xJHDvVAWQahSWsD7vfHPibctKp07V
l4zZAqc9zB0Z52dHLogQyIbv9IvENKtohUG9FfNWHbNRJocAhekqdX7/xS6lr1q1
4Q82aO65KAcZP86qBOwrIy+Sq7Q8z2tiPRnu6jH/ph2seXxjgCTnUCf2wzK3Qq1a
t2kCL/oFmBND4eBjkUf2t7C/fCKZMW1FvkYdD9Stt+U/x9YAeqBpNPVJ5YH8VTSU
t3WFu0wBY1NlYGI2RCZhZfzJ7LdluomnF57ftIdGxczW/2er8R86kVhIHVdwKw5R
pzYpTFeQhxP2bmNxuJF8hJLd6d51XtUHdjLHG+71ZwnOlkaKTTJkUFHJ4IWk1o8Y
dndzq9jgjvPOa8rGGrV8AhVik29TJ6HYoTBBcD3GktM2SobHLUwGVPSj165hZiE/
DoZhZJalqRO81DlfCd68HUdxSVEX+LQy62FDYjlitdCrOvgo3YwhdVUDfhTCkBrr
aQr0qbHQwPkILbLkOpMgiND5slbwdnbHs0y25L02NkWYZhPlwQ/wsI2pZLgxY9cM
tymaNGibfCQqD97VS2dnuKY/JKULysjb5HfOE9oUZ/GETAd77ZegGhxUtwZlLug0
21ZNjAzkIDKQakdRqtXSVfLR+Bv7PODbi9vF1OXlB4kAPwd99YsPU3Hj9XEif+TO
1mGdRkb3SVnz67Md5R1cv6n2mA7HXJG+Lrq94PenUK7y4X9Lg10Rkrk9vXsuZ/3w
Gb6piLMZGWGupi7BQMYy6p2D68qBr0V2+GTxHmaRcBAyPh0YikuSzl3+bFZyI+6I
HHx9OcN1QSMn7omB6MSCudtbrqaSYL0XKT/cIiuvCaTtGbCksACWeLhdur1X7EUS
buGZo4Q+qfITFrqhg+IRW3gZM/nM1ivqR4OBM4sjiF4aV+1+yBRmju+nIoSwPmzR
zpD04LtozuikxoAhO/T5LEN3bwr1jbOvGV9upEFwc7n5pVHhx9SsbQIMbB3rPshI
2igWmYYfvh2q68vgGaVf/afLScAYrJYxjOJjeceRgV0+DjW9I8A3HdMwQTRoCUoI
4ysSo4Sq8fox6zOyKq2ArQZmSmrs5p7Clmhq29bAwHEVQrkKACntYhwcajJAScd1
VWwQt9HaqZK+Qfjqwv3Z1B6pPq4JH+8coyg10Xc2jZ2NbtnsEncbYXxKe1sNs1yR
fTjtiwPFSbD23LUk2Wb5VgmoaZOoTnUsFor57+mqZFOx3Aio59+uWqSgha7CH07F
DJX2sVcsTPmJqd4MX3iOA04KxNRYHsPh7Qf/4uguQm5zvP5xBmJKwbgqeNFqF3J3
pa30k1j/a0SjU5wTk6BynL/wgrpNAOIE9WVM56rU87iPwnCX2Ag7/NgwCyeI/ymX
+LjLOrFfuEf+/1lkOs5hp+q+NWNuPbT3jkrOREnQb0m1dMng4PJz3F0otjElpDin
mbBm6G4Yr8PDnlbZNGjbbVegea9JrVjbUxSQWnJIdUMUdr5JGrKB0ohQLCaAhCzO
ZJIlxUB4Tx9ybG++AAXjeUYNY+wGhrp9ZvrS2xVsg3HDCqRbRNg0LmCcWP/k0ZUN
Qlx2EOR3U4H74SaGS5g5myZZz+/s5LWwzeiqabEUbEUjIK94Y9/Lq/epSCXsl3bK
mRArAN1C3EdzM3zLGrHduTsZh+KfezevoSJAQFEfD6l7rr0zSpGK3oz0pOUjaiQf
Au6IeaLKS3h0JK6yEBxh1F+qiSSmOR/BwAucvr1SG7uTvcduQe7RI29MASNQ4d73
5XEe7lkxwKg8GbbB5tp/KDYg2G1ZjaCSjxuGpn8hjZ7cao0RloOKsV32YR2WSUYh
tHiXVCblT4cLbwV8srilKrUbmFM99MvBn8w7m9nd0C932mWuNVF6zQH3vWQHsPvZ
t9cRkvtWh7nlKDwF/QCPgG8ADWzzNsVISClCOAWJmBGSWt377IGjYuWNQbwbwc1V
dAj7DhB66+GXUhWDgduqVQRoHPfs54OBLz7SUzeWX1EhF1SaUtVhpicycJY5haqw
N1d3KNEWIMhUT8hqfCzusuTbFCtcJMrB3TIe0Jzlx6MNhEM3XkxRPHwUP3obM+xX
si2WzPZX1bL/xfWmyFRezAcnTfrIb/Cs23ZtgOhwRq9nbbBHi6RZHyR6EZZC7bIs
0TaNwT4qfuGOuacswaRCsALWvNVHy5bdreSrG8wMDlgX1VVXU2TeCtrAsWeShCTw
159ICngZPyj0X6IFhOUNgvBA1M2K6Loj+Kwp/UnKC6GTDqfackFNaUNqBdd1+QPc
H6uI+04qtoCiVYoTJl/nDMLAPz1tadfsa4YCVnTzUHrOP6PDMHbMX2mHR3x6uoi+
72pYREVdDfENs2cbtulYsIGZVKR56f4qzWeAfPnX4kWoyQqQ7QMrUfYwbY31gKug
u1l2nLvmwNkaZC03PfsxaKfwnkkC8DQTqbqaASIQe8x51frovTGl1aWYqkOzH7eo
4mthRywbbnS/JmWdYxrHMqsmlsj02vYM+leOGDvOLhCFJs7hbXjFJyoCT8yosOOr
AfNuprarb1zbHyt+V4qkliwzdU0zwtXb3/IRKUVWPal4lFy+OW7WLH66fNfPlBTi
yUvaJptc2LhgpiU8z08CGir74of1SFvNAj5Lo3LQdrcZDuINjRYQwIDWv1g7nr++
8BecDQSRij+II3igeg58K8vSmxY3QcK1/oBZYSIkJpbatsSG01CsNdteclhQU2sm
vWbeICERoiDGIHgi9P+inm3i3vGCNp1MFnh+I47jRXazMU0JmssIgG1cv7+petPG
cEZ+xGuCF6D0d8XGtlhZbB2thxLE9sHYrZVFcQdZvIg0n4/S/YbbJ1xRCA1mGozn
CLaR/wj0BY72qCiBKvMuz0BIAgM3RAEYfha/nE1DJsCM0tBHTTchDRLsGq3BMQQw
zrEnEj9nRcnHp6a1M8jb3jEcFbF3XAuUEAUX+5lMy/khMO3PPrrGjdnwv+B5XyjW
1obBOm19aZOyId0BCpUqG3mSoFN+PyCWXOJteIIT+mLuQfX4+hG/OpcGLnlTWzjC
jtAN0X47DX7vztVYCOSvzy9rwOTMVjJRpUqmPz53zSklrBY3N0yjF+GAuVllGx/E
eJuG3l67n5Blgy98akgvT8MiF/CGUtH96LTqv0dxqJzjixVj7iKkdvGvw4okoADI
4bo3v5raUUyJ3ddxF6mon/Yw8tukB8hf06vhS5ROG2iFLXlXKLtYeZ3KhxW83VVd
6O2W8LB5Br7+LDn+BtpCIp75h9J3xqaUMrVhacl91VZ2tc39xMlA55yzfxm9uNOq
5ToYLz61BbljCBMTTx+RUI7/o/1m40qip2vv/xQ55DIvZJxsXvNfLKk3lO/xyDhy
n9oCmuxvhHRE60IKgf1UgHCmv5AyRZyb9yzkKRGWZt4bKWnvIgOJbl4Mwprph3dU
M5zPkCKAEq+3ptgSLyt310fW4X7J3jjfVmXQ55Kws8SS+NoMjtOyxwxDimT3RF7T
p3yEv5XSNVqQALlAe02MrKMXaFA8xnOpQ8u4WDNMNtCUIfL9i7y5bdMPSdKWfTif
I+kNt1JDroSKQdkVJH1lkxPeK2ZXZkz7odhKZr/ybh3hJ+Y3JoHWcaBh3FosBEFJ
XgNtf+NHSB1eTFS3Wwua4ucbf3tJAAzYttD4q6zDRBMnjAuoW6rOyJzT/PVTWhR8
0VK3FaZQkOEYeJqASHBzivd1earEbfZzYzr+KZXfMqIGnh1MNZ1dSb1QkHLZ66ha
qFTRH7R/9Ie5+SFy4UQwG1N1NOl/60EHIaenr++Kc3RU7wDWETvqv9cOSA0j/KB2
vpq76q/naKD7yeTQV1Ca8yxtbGT7RsvN2Fzxs9scSbo7Z7r8oTeNz75viNFO58wn
DGfez6xKXBecUdde8T+b9mHfZoFJrNTZKKMAn8Tl2ZUg5JCxLjAomv5ROWIFMMGQ
o0ONRqTgaekPRLU9t7Broh+xGMMT2v9jHcj5fx9S/0eoVDJKONx0TUt/uo9YenQK
Kuxl0sN1pg1Oix9Au7fz05d6/Pf+EBgwpw3dbEr+hZ2IVeNeddiG/aSotj932IDj
Ff3DsgbRQ+WaRxSoHqv3EcVBmEiquVQmrVyBCQLEG/pN+RnUk+M8PU5MvJU0Zycr
0Sqvi3Tw11MqgRlEUw3lHI39/DlxlwKVT53FVSrKaOzSdYYUdkZbaObBHRIYA1As
dH/gI3tAhshKeBW6Rt2u5zKCz2+YM43qsIm5ZX63XUnimZo6uAMCVZx/2s31amZG
3Ui3+IIj81o4I1OvHIOfnD/uxxT8mJxfZOfrVSJ+SEtvYCv2LyMvJZUx/nGGqod6
o0wqK1DidqVy8z5rjoYtuD/WSisq+Kyj2ToXCbUMSePixqbmv1XzhBd8d+ti9rak
I43YLNofpquOnaQNf/CjjnLFtP3y0BmMsNugvDjSc4MS5omVms14cO3rnK70/D0l
m8KE0XV2CW/hs8fcby8bzmx7czmHcNE3Ar/e9X6dyedPCV2iXB6HeRgwaGpPucjX
t2YfgTyfmjHwneBjCaNAce33uzSq7FRShcVMfsODs+3uh4HnYzefgoHaUisOmb07
/FzKQ4XddyVjqRHZH8KcUyPl0QN9sElln7RNmemFZtcnA3rqlR/GhC2MLGJNG7tt
6pi3WK54JF7D0/50CNKXd/Tp1PN8tNDSmF8zHOFaw7acqB0nWKyOHSvaG3X0FQd/
sq+bcsLW2NorOvT2mnqgEMU4Bmv1+GbJmzW1YWfxM1Qnw9UWj/ANoHboGUVJP15h
vxY8pcTSFWRgxjG/AGMK/yVhq3M5LShHlEi77b/B84NY/Z6QhlNHBfyrsiwPTXHP
WPPwbdHJyuk9mELaCtObhuNZykdQMNb8rimcy4y9hbXQqSP8bo4tN18bLLgCsv+/
M7bQcjU1Upc5ttlrTmbNJmVm3/mu3q9vl0RFdP559fr8q0w3kHpG96vJbaGTTK3S
BRCYVD0C/nv2LZwgojnMYtrDKoHSqgpdstn4+/F0Clw8Pbm+NJL4iTEsS08FNbDT
lYZ6AjbYfES6RaKuJd2nHKKgEiVBaUScYD18IRIQGa++VFyKo4S6awY/JygHbKHN
k44WPfgVi1dGztqK/+Zwr/+OEmH0C07l7rt69AORICgR5EA/e4JUe3/PYFxZyDlh
JZyaCKIvpT0UKv+XkfgL+9oZyRqHEC9b+CnFYBiXs8nfB0Kz2JwhHrX4zByYhTJ1
GpD0iX1x7BFeQp/TcaV4cgLVUl4j6TLfoYmoBTJjeQfLQ9qsv6DDVMghmP8HeZHR
Y3I1PcYgQTRONaBXAR8VCloR1A5lnUBU5Ii84xdSZP1cVWN29XXFfockdzibsdb9
UhmcCh6JS/99Sh1YlrTmOcvXGFpPalIdOFqRQx46W78eZBvt7yF4+NjDDyKdcJcK
dRXgpvgyOW/yXo0WipOXqmuJrCFSaUKBQLCdOblVauHmWLm9i/LHtzUc6f6b59JG
3wKFD9lYhPBCxd/yp3bVStQ6/ULoRJLkLomq/7KGw7SfqDHtvQ9o+SuaNXoZHn9j
P9O8hnOYht/jbsKoOfroMucFs+aM5qh4TQ9/Be90LsJ60NtfPMUu4JslJTcMvLhj
Yv5dFEgllZV3oZZMpZcRbWufcOqSyv79AqDF+MoJRHMSdZp6/kBybA030aCtjCPr
b5q9VgjI9DuoeYq4XZ+z84sZsL0ehq56g+zezQ3l9fWEoPIBIfjAg2VYorjsPxGl
CWyNt921JtyIKjnCiLujDZ48+ZQ09kgRIkQ5gT5/UnvGVhW9+MgjlTzrT3P47WiZ
aN2EJuihZ1V7krDxTLicsNs4+VK+Mh85b4xEyhgLlnmqhBFHmEr4Ef/gX+/t3iwa
of5RUY42IzKZhamBmIu4eIZ4NF65RZ0Mh1ReHzu2jrdi1hNGf4/x0Su9UNLxJ3Wt
dfCyJMRYlAQMpL+dAmo7rJYSWCJLqIvh/PiYpqG30X0aozpHN6LU8niNa/c4ItAn
iwnYV2SjUTIXYJln/jDgCsRS3AAYeh/cYgvavj+pbQFzfoyqxEASZ5fOrKSSeGrd
+nIdcaW6kDkRg0SyKdOu7JWrj8DDnCpCOaAz1DxayBg3V8ZvNSZWE28DMBfsK8dD
eBlfa8FjopVid/OCanB8MK0i/BKQepfbIODMse0DyIlC6/ZVg3zIF8AYXPSPEv3L
5l38GYhCfjSzhvo1mkYJ9MsSYTdXgStDWpDwDrpL+mFg8UK6v+eX1W6WDWkaQIcN
6FrCZGnBUp2uG2ZAmUWKmuJEiYCIGNXh2VeiVt5TDtJtcnVPyfWclFNGsyGTMZtB
ufPNjck93Fx5j1JFn8Equ9I1abb0V6qBUuWobmlofrKaTjVPobvCJWOClKONPdgY
u+r3TmVVKDd1a6UK1cIlTRf5Amt17TF1AB+aPSHb3lcRqrc8nhr5dcNZgkoWgLyF
HbUCY+KJjCNpT31lnubkM6pC4jpgyffABuDN5Uq8aC772bWwqLiF8rMwKtiFoc/9
UzL+FkBm1twLmJqxzx3L+6Bhru2hcgjcpPZZvbuLv+CMOXveZ4PwlG6cubbY5qeg
IX6oJI48/ETo1TID22vSlcjfz3UVEh2iGpXNin4Khmm2GgQ/28WOOpK1i/id3CA6
pnr8io9mDseqjPzE8o/239sXu4Bm2DDytCX0UlN6Pj6V8JC+W66xfRnax0Ic/jQh
QxHTxnlz94y6MiDiKGkxKWvPmu1sPstI2G5z4IfEX4OE7tyA97A+VEwParHouOKs
XEBU3bQywcHpyouHJEoaRP36cZqEbx6vyI49/RicDMkL0mQFx7hs4zcEFM36/n0z
P/PFmRocF2moXLDu68HCZ0bwcNIsHmBZgh1XS85NwzcgLepqcB0GQHOh9qwa5IUm
zUZOnF9nYEO3ubuGGZ4GWugtCBCo6Ve/VEihnPVeUbuvaDeG/k5Cm7JiiEoi/VQs
d18QbI9Wf4Si3El0unTEG5JrehxpMhNww5I+FsR0tZLsJudSaq9iT+Bp79/cSQOl
CAOqj2L1J3G5URI1sJk7PxOia/kQ5CijlF+o3pZYtbaPFB/qs/4I2XxnDPIuzjrk
/sla5fXNbRDjSMGIhdpUMxX5BXAiH7F/JXeKamwU/1Agr3d27srbfzyTWW21sZYL
Rap/cOwalJX336xNIn7A2DO/3lpg6/ubfA8qM+A4FM0E2aPi9SlvrdPpGXvZeqId
GwC9zO+S4jwyAaCLz5XcvHygHB528QIq4KqbCYHbjEhRksBsf0ZUbwvIIlZusWXo
cSUl/L4+LxPm+0ODC6n1Od7+vtLd1JW5PvLzE5RrXURevWVfPrF2JqwaFMaCga8J
MjSe+NVF+m35uyiNtzdeV4CF6ae2uJxq7rbn1pJA+oPFNI21gLDVTkvIFBd7W9YD
GdA6GuVPFKZ1p1NRqMlOFMbHWIxG1VMdMZ4UXwcYf89WmEvyT32j9k2r9L/KUhhf
scI0gv4zH3jkmgEGllIBa6jgwHQzsaStmpoCb5KAiCGPVV4gk8j4wxeGGoD6FjDT
udh/RgTdjnO3c6bzuOwIoInYUAbmq1Vyc1m/9T+68SiltOSYBQbcnN6MV4BWPGNW
qZfqdpYJkY3nhkP3Yoh+Xq/Av8JJSBqbEtRP/XIbazu8W2kMrpD3eN4uEF4+uf93
p0azCn/V0RVIsIrY64fvKlEDVsdHrTrBHR68Xdjr/9U+dk7hED6OCeatX6INDV8U
ZVbZIan2xQlMDMXE1UGE09y+5hFHipMru7yVWG70JGWsNH2hTilmo2VbmtrD96mw
JAsPFSE0DvE5Sd2O45yeFBrupBGXv2EiRSSie0cd4F5qkHPtttvPQqZ7884WXg18
Jt4F06cRsqQHTTYrHS0ZjTLVlt+UKcObBUtbRL1hqNkOG1DM715Bga1BTuoE82Za
HJZEitOvWUtfVyB8kMELyIRd1mNcwXffX6XgCgbJWmJXuDVbQgfWjRtVw4VlW4WK
XvkzGcJFq8MTVJnqD9BSytqx27EZ+PRxLlO+ATqafVd7lpZd7qe0HtEdbdbNrA3j
IdwTyWYh/hzGgnCdxCQKn4ULHx+mM4b8CDyckkuCKcnjQ5RqWqpgrYbdXRDPIPpT
YgLwh165TpmFVLgYknOdwjuy9eN4oaCU6oBCRLFkMHGoTqDnDxKTFyOy1plJ7K6r
0mD/uh8Hk+ku/OsSV1ojDPKcsqa4in684AHdcpl0KVxihh+bf0rQlcy7kp/fTQFS
rJNXwmW6RRlKcDrTRFvRvdFCHuNPaTFuPBsG1fKtuaaEhmU2eKrBxNsSATOkWTDn
7KzfoboCHFJrcNO/PdTdTMMS12hBw1I2ZoXxFHi+tyuqT6q3GwK+ONgyqGV8s/Lx
AlHzu2oYIbONdnpznKpeNjJ48dvuarS1zXl/3LvPh0LLV8GFCZmskikyFI95XnmD
n800Yuv/0a594AG1tYfV50JiLLai+9WHJ4HBsAOC7xnsmi2toJVtkynNprT01tXL
4Uulg3YoUfbZs6Hqd3QYLBc4Q8Ws5sQcXno/7gi6lM85yTC3xmdeJzDRsAkRiWI/
kyuiwLhXya4tut/k4v1qihP1LczS6MLN5Th/SXLThM6yHLDLqOVHfJwAhc9Xv89I
tdhPgtN5S5jUFvFNWt93EKoyNCfPWzDCvMEF8Q6I+WqYL35dqPY+wDXFDnRQPU0y
1mUoFnr5i8GggwTAgvnTeWmjia85sGrcMsRIX/sSXMla/2Ij/YIfC/GxOB2Bhnd8
xtDyJj9h5mpLTxPomGTHvb8vFKt8Xzg9GQUyhIFgfa4y/LXkepsQ/55pX1MZXuci
voxGnx9uRT/j7SWGA1STEe3Ys1VTMEbIOGiOLScFA09lvMU5BuPi8iEHqgvpU5Fz
YHvD90pv0Ml7e67o7+kNlbQsD9snZsBfGQacJIw39DIDl3B33zgDBCIz8k8Fxry5
GRKQTvGXXe7+AEY53t2OnKQ9mSpnK9TdPGr2K9pyw0alk5d9F0URVVdjGUsvmPXk
p369iwVqZdgG292bjhlLQRo3BcKxsq7+PbRrnsH+DjrUdqAX/z40wXdOamqcuRcL
i150sg26mJVLKEeLGM0D6KCWMLAVdMwUqUY48ltxXDMRG1HSeGxNPus6HRloBo0A
X9c0E7voRZlu3vQcbXknTc+v11azAVXv4aiF9ilFizSZcbjJ6IV45zCrgBKQaufz
4e979tfmfLAu54DZxLKfi+6EZ0yDgsOclmb5MQnvWowIAj8aAqKMCFkwg53s1Wfi
uvD0/VJJCfh1NS5nJrDMS5eExnqKfv5rPS/GGkvwYJz9Vu2XkI4ZXoZy4R7xIxOG
KcOghbkpxAxU0b2f9cFOU64CRpQZjKPknKj4wQ697/ctOJTZdEqMbwWEy+FjPk46
MlwnQAwoKFmh4BSqE3KEfeuK0CtAPtcweNqovRabQ6t//adPE6FR5z7WYXB+frBN
xwn7wqchnblhP+HQVSrP6tMN5evanRthgkfCnVVdEJ7I8i6kyJG1DisfH8iPwH52
0oVa248fkkkiwPEvish0DXItsqGfJURP+1+SulUlB/stUY/Ej6krwuBVJ7aJ9cW6
llMHwflCDut6pRvn7ygZolAudT6XbLHRhDwBDQahkjmXc29ya4H8mhcKDxzqFuBu
W5IHHZgwGSQY86qyLeoBLCHg30GiygMIzcHyoCqs9kKOcrDWWRBxgtINvpX+kDxh
zRJIdNhtbOINRZhJi0dEj4ukd8bqid5mGgA2jTBRlbo6otk1v59P2nT3aabx2pCc
c4N5TCimg54fc7itC6qx2RLagz4or/j5QUZEnGJOcHzbcSsa5BIZ8/YF6Mz0vCxj
ompb+NJVBWoM673Kh1EEzNcu3VTEs2UVGy/7dloOVbNwT5Lf8qgTG33xVv+kPk6P
AcYFHamEIFtLu1s1U5kqYhfidEYgCAZaQq72X1FrBytX1aBOEI11d+ZBaY301SzR
q9ScyQNF5ykJ3iVLfawFdwvqHk8nJiqRLrpBYzjqp4zp4eiEqleZeoP/3Uf5RkGe
sB5rOrr/HOEyEWcDmdzhM5eF2PyRj+yRMNH6IINHV5OecqtwnLejQ4J7tgERgaYj
G4Gkgd44BYYIfuvA4Q9+gXUwKFohhEerkR5gPUL0aTNTVIQZpYvtCUrNZ8T4eHqB
h7JtSmHUsAD5beQqyvHLsLAhgLgiDpsJSXuYsIDC/2EUTb+j7unipBP/GsB3FC7m
2sWsSAhADbjtFUZ2q1gVehXaInENDDCfeumFqyzXIBFgsQAu2AYQVlqDP4pLt4NA
p6+FXY4ZsFFQQm8jbbsk1Heq6Kz9k/HXjRA72lGlD62Mm0ZrMLGHJwVmbPQp03uw
H8sIXsw5C8M1dcHnqSBgPbSbn12w1RuPer2gaajFgcbI0BNQNEHoh5pHA4bCEUtI
Z0fb2Nu4g+lSuHUbBeo/geB7CrB61g0cXB2nmvUn1MVaH+vP+hKjhl0+i+H0rRBr
rGBibDMcT1zMZUkedLgfi7SSQIO2kNx9HVZARkVSFzY8MMvGyZdDe8vV0U48TLbz
Fv0cwE2sdnmipsrM8pRaIJFuHYxQlQNtlOBhvYzoAOGvRw40dtORTiHfbguLS4ba
tBqzQTnT5WjGFAKBDuTjA/tW5Tifct5lOYKxYEpt7H0rSuhDK+2ND+ThKvHwKzlz
lP1/jDq3ivPw8SzdfoEsN2qrZjFqDJ7uPia+lGmpsAyxQ1vVCTX4bPsnduhgcloe
I8FT0m4/4rcisgAZMOnCJjZgkvpBrSIsiyoiHKMn0h/v40AzAdBfKaDVFHRF2Cbo
vVC4tH4HMfFCzxGvYB/8KPY2kvgwQAIh2q2/giii99k8p7c0kjscfA2mjTLgdIbT
7UWnf1aN0NupBFqXaWWNL+VZFMdRSPK+CBRCEIDFyIt+RAuXqu7tff6zB1o5XRvN
9Hj8j6PgcZH8jKpgOEtzxCvASxv/sUoJbVAbSeun6oCkq+AOAXfSPmgS40IxUaq2
9CiJPBW1TQyd3vXzH+rAMKtSl24L7yK4hCDdCLhykl1iybDEAjlLLeDCffsfb5an
d+w9uR7VkyqojTLLpQw1xqIJHykPdqTdEdngAgyyQY7T/OFYzwFAccx8VLQuwhmA
agNhefDJvY90+bsuiUx0vhPA3rM4CnHt/V/kuk2xoZJmnCx5W7TxsvUddTKNwmz/
Rf+D5PxNk20TG/4tfFRqKTsWu+u0E/I8m8QhwNw/OZR4iValScn7+tqi29PI7+E3
A1q2tp8FeTvpQm70ZvRETVNblMXLdF/weqb+tTwZzZvl/YoCIRPEIIH7hCgg0M8w
cPpjqoaOwc0o+gEIxx8suwvEY5VEPsB+5Wwvta3HxyowjOIhpijwHziPX5gA7jui
Bf3PykZkJ3wFRcujFd0wqfia4GL4DpoCchtOzt2of75++PSi+/IfPyoIoiNFKRpq
1y3JvBwXr1scU27op3gORR0aHZ+2qV6c9lpy5eHVPvSnFWH/PxmfubTOAg+LC0VS
KOe+ZocPr0YPJnHAB8Epnyvfhnt9RZ29k+vjI1FmsU2F3wS6vBdRyj9AOc/3Ltxs
ExzGaWjMOL2eQUIafNg+Qs/0B+dIXlm3Lp2CWpZeMWkn4zYUDtX4SodxKd+/stm6
XjUPZLNQvbO1f9z3dXJzcVmR32JTipoTxMoGddCM/vpEpCBa+HxGNmv/xXPmP9VN
6RosgBO7DMquR0zFbjiaptm9xPDsx6vZ1Hfj13ZfxFo423Yrnh3Lzy//JA/jqeBF
IX6auB6/z5TMuq0FYWdlrteBg9+jmo4lOeP6IlCXdLgHxA0QQQmiBgV5vCXqL4ss
YVCfFAlAEUL1//iNpktmsVNgn0UB4YBAQHSCIG/eD3LF3O/Tw20mT1jr2rktolss
RnKQWXAnY5yCmm91HbYPNdNv4fHFyHXjxYXHkfLOP63NABPwQCGJ0kP1aRvtNuBJ
nBbTI8kMx6eBviTZWNO/cBDWPqojXHQOdaOFf1yXaVsqcjJRcPPPlSgluHcNJShY
e/f/QvuLqFwIFvBDFMOpvB4D1VYSCSOb6CrFyNx3OtjMkLKsiISTiiemEgcWB0b4
ktbVJKMVyZF138laFy9WZDaxdzhYuXFfneL1myfLY5oy7RG6d6ptPt8y3Mfbglvr
1yPAfF3a57ivXvMk/vlRHtNqxsgixqzM+kai7nZ/YXkUDTlpKQsV/omp/th0i9NR
ZcAdjT1nDH9m2jcr3Jr5JgtIU+iM43WtQlDugfNNhlv+aFB3LtGbnK6juwfPWuWa
wc2wDYRaKyPE1GIHf/VCHKrodQTn8lKGzzX68I22vmLPnvE6aJnWvYjAtUqMhwXa
fS7I67JJ9cb3tYFrXPyL01yf7b1yiirW3lsIlvFenPoQ2xXS41w48HQgqx3ejVHv
POU2w7oLdgHux+f5NcNoqz9M7Buz6jl/JsaYGCjz/WEmArKXDgOIFgGlfr4jLRvw
pnsJseoRXkN9khUfWPrj66QlTetpOu2HU5zPBlIixKazYnjk2z9AvfX2+JF2f2p/
PCNF86bA8Kf7jwsfSw7+7BCYYXSI1eipdgbxftQGrvjCRgdbK4HxcoZ3wy5bRtR5
AQSO3PiGBCSNkdqZHKVCTHctx/pqYKlt0Hg7yyLUWCqYXc0EFxP5NgEiAMRT3Z1l
8JVL1uUuoEaD0BlLzNSpXaVRsoiskZGjsNAjqf0J7HLxmJa4AE33rWmnhWnuFKkM
bvwuDOJ0zhVw+M7dyfZZGPoL66FQtMwQilOY81I7rAgq5WLxlwptXv+F45POUOLk
kBAJ8Qg5GwEs53uCWtEk1XySoWvkblfWcGmEKIZVqPWTgN7wpPHwwZDQPPLhueUU
TGFoaCnAB67MPBCpFBDS5cMfGyXFSZXeaoUxCCLOlZlzOWPLhoGzqlinHtYx1Tkw
hBB8uVk/rJIFiE3M1Ddq+w03sRHBxdsYnA4QwXGK89eZNV0IFpwJYjuxvyzFc5tp
4lQZEC06dvDA9cQKkbig8NeyLH07MTmIlvY9oUlpID2KNoxkt9ZI15FXy2zpHKHl
Haj8tFX7t/SIO1jvW2R4CeR2s/ISLqqcQ70hOuq9CxRgu2p6MZXaW2PggyrWX0Q+
9e91+/ZGocy0o1en5Mi7C2IBnkoQm22E0jdTubN6D9QZSPc/GZrSvR7Fi+PTEJpu
dxrstkComsOPHZLYAARSGnr5YUyDXq/23mnsvr9Ko+x0J4gx8DZAKaNES+MlZyNj
ZqrB7SxY/QvCGDCE2B4mTHuzjF62JhrSN3+jAyvpxMauu2aSeJHsGqFHJDqUUtDA
j54q3c09+Vn+Q4MLdDhY/byBvu7th5A5DjYA5kPo73rdazFcA1gV39QJKgVai2oW
GLIKd9R6/1xLJGmdRRq+uat5NF39MHRWgivaYUeTeiX3unp6TFwtKM290LjeWU8h
b2UsBng+BYBpnjY7H65IY2YPSTNsixauK+uiBnHkWVDMzCM7m2G1yokIz7LdHztS
420AuQL8cvaj8aMwOmKHlq5d0WG2hKeWHpAuSztbrjOnF3izgRrrXXNjmFoZ5Tbo
WjF+/C1re0GfJKlaZtezthvuZ5LjMB/lWE1um29/cNFTcdK9HPYKqFw7u48FBT0r
pxdr//jtO5XlwNdfKEa0kJnd+9bla66MrtUsWUjio/8rwQEo4waBQwg4rYXvV7YB
biDfbw3z8KkHe4Xdxr1K2zUSZLJPMG2NzUDCATPtfR1VVbqzaIvj6I0cKZ71ceK3
4HpXmsmr1cGiFruA9qEirRRkJ9BsjgiJDY/N0UJIHA1K+1lg4cyW860rGLyUnlkw
xJeNbc8K0qA0UtH4zIbuJpoG/Rul9Eld+2Tz2BwRlG6jcIu7ApG5syAOyARL78ZZ
lLa6zo91SOAsUzaEeGWbq0F4kpMrAAAsPS0et6B8PSnOWlijfspcFKOUbavEovuQ
h4mWvfvXga0xW67VsYmpfmGN54VTijPFh1saIaTda6bmyPslYjuw/URlgcEnR2Ie
hRGN0LaB0jECHTy1FH4mQ8RO+32IiZdHchJ+eZgOOZC32J8dSQnCxhqH9UhQ1Zpd
SUKTxj4tpkW0NFJrrSP/Aag1Pqt0WaDWUkkhiODM/STC05TfSner3hJy00rYITkH
cqyJhi+Nmp8HKLDiKwIjlysDDaGIYL/VF3QQrTJ3Pq3+UFxdZff9B5Ixht/xDAf6
0wB/SQT2n3R/Mgu0KNIP3uqqdLzrb0RD91PcCuEa1Q6Zt3pHRhBgYN1ZmrWiIuv/
atl3S+CiFcu+595+nrPT3kvcwvE6YcINaRRHdq0j/Z8hBvvW6iwpN53ZYZeeoabY
sgoe/GMb/d6lMfDhimYw5MwBM70t8BSmnt6bY3/iROUv0BIiPo3a8cryzyNPplnx
SCMDROSD9Rv6T3LJnu0l/zOW81tKS99eXNOeTRaYFklNnKOBCHwq1yd8oSTmyo+r
tMBbLyDCDG1N9cwVVVxgK+adRsVbBxLdsqLEoY/4QssEmNGgE5tHuIAi9j6O21sp
kAffb2F4hZPyVtJCfG2NCsXtFV5XxOP3QEGtNpcrXdvdYkfRPDVLyZ46J/1qXyCT
bzysQxUrTvAsNaihFlcYVWQGLjQiLn3sGVOwRNhtD0Wks5yt5lOE0t6cCOIONhim
Z5gleCpjmMIdYEUKSaOb6ZRgyDq89g955bBwCQdk/pSpVHKwDgXdCQpbMld+6gOg
/TDxcwp6O6GzlZ8ZpcbiURUyO6PF7f4lPLeq63FHiIV5yiUKzARGSIZKWHHDhKfl
6dioClvUWIeTQBZZA3MeeINWlzubs5MJMAozRckkBuRtNspmmdETriDCkMnfkp8Z
XDIoPxDHeZfZ6AvM7csCpyus7HyMUJtrXbcGdb01SNQ0T0V9rRT7pb/hZYw2px3g
d4vMojDRrb3+7aa1CpVjcjWwGFgxVw9NOZC5NnrAZ0vSzB399XgTltaCN9rLJAlK
X/GmQ/MldFwza9smCFr2AmYFPR6wJoJfrtm8+8cJPC9FPqlGH5clsr7Zpb2OOX02
JQKg+9plxs+QTMK6/b6IeM8PLx1w+7CpCrdS53OMVT/wmv3f6H9t7A701A8jCCUc
stTZs9hDbWQf/1d0kYIOecIPgyeuywfQXHcLmz6C0d+OwwUAZPeh759IUJRz9ApK
fS6xmuLIYqOh3H/6MTOIr1gpjMrRvdg6crK8d3fL1FNGVMyCp13WT4V6fA8BHjnR
6kQhEpXWlsQGOU9Gc2pO3oGgNY+Sb7KjXqQTa59ycPpzJCvFG7Lki/ERqTAGw1FG
s60UHmewymLo2qlbOTPg/USs/Qe0rN8NLK12FTL+Vaxd/XmlQcGaZ7lsiBuFCpqz
yYbzqT1qVFUSesFGkxg3Uo8fb+Uqzra2UnrVeIoSrlyPs7mcA4EbZui8Gd6FQzD1
T2pBxOSFSx59Xvaw0o9oTENI7VCpY6oiJvBU3Kp0KbxDcQu+CgIAuszkbbwt4/gW
ahDBy40a02CQCzqZeq8iWyQDMPBkcJdR9SMlKykVTQGec8H75XD9C4mt4d8NW6+L
+krg/JVGs0K0OSCC/Zkx8FBhWcfnGmwSH4Xzz4OniXRIk++tyToBqParoTqZ0OAB
elaGNItxgCmV8SWRUT0XNWPmIU1F1UKju/g0RZkjwW1fdERqotQTg9EtEjsDe5Zv
p6DB29wVP8nH1m2RImzl/IgojuN8UsdmO4Ay8cP8cKU/EP2FQk8rkcpCtu9cJVva
78EKscCd6bslU0eixqOs+sHgSh5I5dFYK0uezvhB/vewDZEOgUO/VnzVjLoYk8eu
kvD9nvyM9LKu83ibJANcJNV+HI0VGcVm/kwYTophCHq03cM/PWr5DHFzAbNjbAWB
jyfCCtB8eyrYKca44N7A3gY8ZdPoDyv0BE65hmm0/UYP4aqjq83V2mGIiG+vLBDi
dzbq9k2c7VRbFTXoEWkTXZYKu8Zt+bYBXJHcOIcIx0LLcnSKXN5tfcNXRmhFSd7U
naKndIGT4CJO1ySlcOHz0UIPtwkrZn3vQg4vtrx6tCJCrqz8TG/88zsUKtLeQUCp
pc7Oix8gv0Y3J4iX/k3IX29fVfk00B+VxrCkJBpROhF8BhlvqkDe02DKgqbXX1aM
gzp1AWunS7DxCi5VuouGts7peky9ilkjwfMrUXWNaxjMOugx6W5HdcUK7iH27qEw
6zDvp+wuxwPItSUXDk9gaXSzQbx3p/dF5t5U6ME+pgmH6yyGNFoVRCHzoswM90sl
0d4SFofkLS6sjzogxFHaJnWJqMK+VMq3w/IXD+Ki9Dr7lG4BiojBXeao0qQzHiQ/
wkeVxnwWz+BwWVFS5xibb+N4MEokjME7XUoVPxDoeA68mI4QYqsx3Jy8y4Ez4G8q
oyb0n9jCx9NwRRPyS4L1Sv4I3utSovaQAHbQt0JaAoxJNJHtWhi7XSjbaAn9YXX9
LbckGcDWD0u7y1i33nQBQRjkQZEJ7bL9M7fBNfeyv0St6at2+QMslsg6zrcA0mkR
vjKJWU5ycomPSbolFfqu9Wse4UnLLeV4F25fb4sof8SiLHQODe/SbZFi/TQxYtsZ
Si9IeeiXiW26xfHDB0jWDosejVmpwjWC0vAetFXZ/E0vWBhFMemJ16Aqmgkt1mFz
pGClwjZw4UJOIoNqqt+Fn0ZFygzJmfk9BYz7+BqGv+niXecWld5agBlAbQimlCT0
IL/KylkkHahnc3bGfeC47NlTvxJ00EkNT0oRmHTyVcRMQOanLs/wEFXkjc/AYW6R
qFCXWsC/rN2KbUSArZqXQNxiXBFAAYpuG8rFlcSSq493MVkrCgEC33G/mkI3ZNb2
YDmQv3qI6PXFTz/BUXFPJj/VJjZbu/LUox4IEiDfJZmrz50f63LVJZ/8sWkydstb
p6B0n8Wn/F31iBPzYG2tRevjN8Y3Ha3s05rLGKpTkT8Qhav/62DXEE/6HuzM51XL
nWCdYqe6Roa2b9FAbBFKytwJo+8MsTZ2VCctUdHyxPIFkoiY0ZSEu/hVVoD+/Uw6
Xs2pqH4+l5RL7iWBqGBMP7vg0Sqo/5n5Z3Dd3aNJp+YzCrzl23nhJByiyv+Fil4y
8PSD4XJFaFEAmgkJ1gRf8icNCT8ON4YSlNiGmwgZXZGsomAWPKIb6nqgVH7nu8S3
bWjG/MkdjpDQC2Qmo1L0W47JkWyoBu01K/us0WtFyrTylkk3vMnMTEek43MnmWOh
gI4+Bw1/YYEbtB39dTsF8WQFxh5RCCrbK5tsThVIDcPREbg7Cxeb3LtDvK49RfSb
IKU0uYcyeCtRsBNp3kGke8LNC3CcWYa4Rd15aKp/3RgZcsw4cwwUZ17qNF9aLMFy
rWdi4Gdlla25q/6zctIhLVj17fu6l3th+hDqG7rYY6Qb1SoZtYCv63Ga9Jbzct2B
WoEcvUiOjwR1yhIfHA5ZioEN8HW5cqFY0ANQeJ8tVvJT29Y+6Ed6MEjBGLnrhvxL
RfVe3L/GMVJU3GEwknPzUlvlISf58MX/20abUN7ifU1kZ5lTiDnFxqmtXu/JS/Fn
xLmAbFvnXE+bHSGtp3i0FvrIVVVtuXvmtGRstiB36sxPW9owfve0tCxn+pGv96Di
BD6iimnTqer3QP7ppVrD3kW+2VcvmlXiUqvG6wTmE3EZHwHvaVzFSJauffPscmo2
nQyUcy4bdJ4FOUmDloNfzbwxZ+hTxuqNjD3fQ+nAti+Ix1JtmW5DDt6awl8pHpui
E8w3f5CpyBRq/PlpEr4ixfA3juTcQghNAZE3ovYMbzSvNji1s3/Dm2qCAAL9jMs9
/5gjQs4u9lP4VMmXsrlT8qWqB89uImC2ptjEWmiotFDl+mc5bDxQTiD+/78or17q
K06pud4uUU+uIzU9HGUzITT4oy/R7+pXejVRB1G7g1AYP6M14+38+rTld/H2B7Ti
ksQQTyx8FKiJitwKrxczrsYC+lpgiO8lAQHpdbxIRGcJ+1CfOrzetF7uOq5slEeS
XAEoFHPTA5bbw1UycxfbZlJ8G10pHhDKlDtMnE0uef9nbMIuedvcq6jTlnGmGWZK
l1IXy/dMcEqF8KGLZIQQKe3HOUo+zNBmlO+1NtIqvvq+0IxCKw0vtHmyuyFlX2Zd
MSyHjAmscykPv6JrCZeHwBoQGOmIQhhTXPlxK4LgtmbUStEGfLm6NanU9VnbVwxW
OkXeXg7YxIFcQl7Wn+CtmyQHYarK9kBD7Oc1sNfYuVqVxig24mbOffvO91ulnaWH
Guen0lPMiTA0ABRsmWy9YzKce41oZlrBBSNWvSlKqfPbDAmEPHN29K9kdLIaU1Aj
Y6nrhhQzeG5YFFeOu3HXJZ9f+NuHu+cH9z182AbdoTOujhpUf+NawIf7J1s8ZKCP
MCLRUNRJx1bJlDFgiZ8fLpL0vAL//hR/mo+qEqJ+NgaSqyFKEmm5ccmqzfqOLU4q
VwCKtEHe73YrypA63yHWstLGgiRvWay9ZbJSsm2ZVZzTp4mkwGvhNH2ZXT4E6mc4
WgS+5Dsb9gV74iKqePOBZpY79wQmxyMzaCLezGBL8VblLxqeEW6HIX6m8GJfeGSy
70TWr30fpAQZawdqqW09VFgNwiZDsnP8T4ED9XnOthP57gvc4fKDVqL3a6/aWAIp
jEMmCLgrAQC/fc1AG/egq8/H0Rpya6QNyF0nANVV3Y7PW/TtwUTZwaeK+ARYtgL2
BCQO1+fzUtZupsMtFnzRwHv9NbFwJ8Vx92NORhSESLrxgG0FW8bm5fvgl8I+XHK9
M7lBbNqLA9gyyAaCjYD5sEgikWnYiFzAEjKrIcEtPg9/gnJBDYE8SG6NPYFRahz/
nxcMHbmaV6N1MKMXu9u6lV0cEaNkzOnv9SJkRHCHFx9X2Hj3+1woi7Tw7/GUHKPK
8nHHQ8GU+O0jtSeLQ+Ffxf6J2dRazj3SuMtDzXMPZVn+ZghnIvq3oYfl3Xmv0Gbi
6kojFYyCAxxPZaKxM4ZA9EObiQcVWwNQixqOIIWLFCZWDa0+8UZkQMWdwo5LFynA
VoGJ/IOXh7vhym6UQayaSQDBCUTgmy3LPA01JRbVsdyF/Vmnpn57erDRvIGJhqI6
YTqgz9qgWvJwHIouu+TIr7VrgWtp8Lyr8ds4kn+++6KKYbE6OLjFL4MGFlJPNWLI
we7Ql45ko6G+lXDfKQMEzdjPjPhpFbNgDfyaDBaB+e8q4tAppBzCG+k+7cfuM101
m4fJ/sg6aG4XoPtr/5YOyDjnFcOjrm60wff6L0Xma58BBL071Pf54bKPZ3ki5f2f
HmnsHYpjcp6nPRH7DI1+Ngi15CJj+IHtDcdJsYcGaPurWv7zrcAGqKpTQTZT0EDO
r7V2ZCaJj9eqmsvkjczFRmp/9FMK6RE7ThxoYl04PJmtXeU3Cua5dZDEJuqwu0Ps
jwdIwPcls9YeoO/OcSEeXNQ+mnPeqtL9EDnZABNdL1d7T5rPp9L4IFMsHAIsYF75
5a09S1h/dxrL58Ob26gLJ+jwWUHWgy2EJToS36japLdPLtmQFf3C4LqFENoYcCzk
DfAvbKdgkNiSQ3ukM39UJqUxXwiL4kP6lhHN6NA4aUSoZz3Z2DSZECHT9xr3qDdE
E2wjHaAqZ8YhIYSlsxOglo2xx0D9CTg9L0D+pToe7NRb+eCJJXc5z1iuX0Y1yiCS
khVPGQZMhv20Mck5M6WTVMfN8ouXJ+Tg1q+l6mGhczLKXsMBCBMr25KjqgyADn77
zrALjFcmrCSm5CmwHCZUoR47829bXFOXJgXv45s21rhnunpOO+A7p7xpKip25KS1
Mas4uVIaBlRarKJIwcHMU0wm6znY3i7pB0hYmAGlj2A/4gmd6E/u1AwGsxtOCaix
gIKJOR4zrfXvLPhQ8ESRBG4aTAPLUuibLx95XhNVftR5gcLUxdHQsC1WAQFnxhTM
LdfYWoI9Rh9auUiRTwh7Gqn2Vo0wOoHH3aidcBSPVvIJ93EdYD9DQ7R9EmCJyi9I
sAXnt26KpeGpxJ29GuwWtEKX2c+7972Mizawc+MjFE23CUhUcxjSk0ULzIwgIP8Q
UqT3/39kkfOlSy95pfrtWRY0cNonjfFF8go80lcHjKAyRPseG7oq31lTegB3OrGZ
dNgc2oK+LqD3LPWKVXI80nAPulg3+TG07GEwbToxFCoGuGMRm7lT0iAqlSiQhqtx
YMOWeR4U7o6p8ZLQjrBOEA6Lal5OAsCj8hR+EtGOc7O5FkehlFh+4CRGhmKojzaG
zn3UUA9Yi+F57sKHUXDJdSUloT059BMUsR1P14UMT22ERJt5BwHILj4IjjJQnFFg
Jyho2Q8Ek1Ypyif8BEaO2ORHxqZhH9t9Akcd9CPx/3IV9XM8gjXhrgNAWWqnNiN3
NCAcLgRfSzQVKJeBwh9d1UbOzmfyBhfVWI6Y7XUCYga/plA0w184DhMhRbieERBs
wrVioplgDhKGWec7dZAyAsi/8+NmxqX+mUFwCpGSUKSgzZKyDAW2QIEKyA7/wGBz
GlGwjiTqF5AXpKqDGdpRAntdVONeyJb0LYaoUbsTF5uOtPRZdw/pna82srm9xk72
Eto8ope6PGUEugNSmw/sC0cE6PrUKE8ltt3G1nPjmbvk5C+kJtx2OawgLnMuCoQy
UoZ9/7a6ohRTyl40vlDY83LoogLPql3ctlS7qgo1nVT8Gax6qX46WOmZBfVBGIXd
+wIoZKC2nv56xMfHvK+S/Tbx5xcOBOxRiZdraOK0EkyO0c05WwrfSX9zoa1gFflk
MlDYDQSS3QMXc2Z22TILtGvgGGDpZXmTB05GyaKR1DTRCZXjw7YmhfkU0BhX7kLn
Vo80WWNsp0xrc5BDrukuKUqQT2ZdeWFOTZ4eWscuLtKkS5lBlFRh3vZIgv/hkT5R
iA9ndQ9LXlM3q4HXNRwg21gI8ijR/Bpbu+VGip7AfSfNK2GmkaxZ7EctSSNN1jVO
fRl8qUP+gcE1DGH7oZ1ESsheJiufFu967U4Xvf3YIr2B6bpoLm2VxNP4UpheXppW
LIpnL4WxemQCYg85rXrkJ1DhEiaftLnjmzWPFhymY3O7pZmO2P5g3rHercVD3s6T
PWUntuKtJmtXdJRe7Re8UsguOFG6hraUfw+3qU2d/eFkGubD4/mIQn+ISp0Z1we5
BTYQ2Zag+NVFPmy4rnuQsnHG4a5gpxs8lMCI3wyxBUABGYZYKz2eS8j6c0EG8CWh
ukMWywD156c5zNKRQedasx1gxesoVUjpt9FOhMx5kBNvE1bT5DVvYXTEubNiqGwV
+gEoxejgoehI3PCrkYaVTqHCl6iHtS8xB/G658AbVEOjKbX7o4r0sQPVLvwFcW3y
rK9hJt7tE+NGknSzqWuSdqfgV7hvbtVrygp0PwdqKNms/V6A3cbNs1kV5iDVapaf
7tea9ABCfVhCXZxUGgUdRbB8e2XZZkgZcGGjqJOdSRPkjdohx5oFJqt5hyTJ43qH
zXYbvyrwPOPeVWL8ZqsBeqqnzbqv2Sp6imMBpf6KG0h7sM1JNnRbpGxb4Lor+3Qk
zEGq+ep2JVejBtCQki0f5/T6bqw1WUkm++PLz7T1Jjdqs6S+sPgQ4XH8x0v8EuPn
lFnKsd4PPW3DjGgLaatQDOyPEh7JH/YG5XcL8H42ApkRcR1m+wEOiJ5UcFNP4ieG
qW/ZIWh2/sNsuoQP8KZ+1EYOoVbqI5DPS2ToKrqUazihLpt7LTYXiFnN2as5pp+T
NAEsYfDZFcze6lqdkZr6mvn0EqgLxk8X+TT6fUPPvghoJlB9ygvLsQX9K7ZuJf2i
cVBg9GDxKjvxTB+CJqQx4X/IOsuGgfJdLDgeWfaykoIgxGGmLKm7nRlapIsJE3KQ
IzEh20Y73Da5uKfLXXzxATGvTlp7L0NJAlrr1fBep3kfUJ00F6HaVghIDU45acMo
0Ci1SENNcf5nu3EDBDIsbMHCDyLRGBOf3c+sbmxtSTfFnXUD4CDO2gSi0Oh5daP7
LzD6V8cfTH9yso96xWk2/0fCuyINOlaxmo/mzXdkEafMWgIYswjQrF+0oliT9uQz
JT4SywEi0uHPmWtmtfBmisaRaTcV6wWH4qsWiwrDQjpbNnLJwT1nQnuyiYuhh1JO
ir44Qp4SzuD+WvjJDSS0ac0kwxrCZJazF1GN6+UKf5rzWOYayMksXNMpSanoq+Dy
tjVO78vhII57mgDAjPteeZRr4DoQl8DcY3UEVyMBaP3cUh1e27FqN1RTtVQEnCVK
n3WYZZpf1tRsV92tJzrGYt4ZpDxdE6RqvTUR1AZ2BmRaZs5tyCh6LxyT9K9+yZxr
7ffEwr03sfdh4muCQb3LfU6PK9Z91fCa8OjkN7lVVOfc+hloaPmpO9sYPQqbO8f9
s2hivIazYipU7yjSiEFgK1SdMlKKnVP70SFyy/IXGEFD9cXXEfJxGCV4XBIHKsvd
uqm+uIiQey9V3OfQcNmCnCL2WzSt15E97yoxxQJcsEy9NJSlaTWc+6eyYgYzsun3
iOHBaP44nVKDLEYC9sVeQO2WMtNdJxktt4flRXfroHCRUTaEJ9xLyE1ssizRuTnt
THxFu5k8sY0oRVtSkfayfxT6kyYaevPtQtUdliyBoar8HjdggheepLzp1+J4QI8G
8f1bBJsaKRmFo42IP4eBgmLmXMXMctd4mV5OeGJ8RW0yxhg98Shc25tFb/1aPOSb
IH5uuL5aLdnH8F2NwkUHFVY8MjAzeDu24xhEh9XnoXqY+GY1wEBdHM1LNfqjIcBA
BKznv5WgNrDuZOKgbNAap1OoUHxyoCnubf18tnnKUfpK5ebyBHmNi5aCuKp3Ts90
qegfAAulzNGzl/xPX06BnGp6i0YwZPFa/teGjRi1m/D1JZfd3dL/DGIfVzwckExG
29DvDADj+yEl28iYruOk0tKdAQS+KwbNm7JJ9DU8R7hYe4AFEsFrOW+/x/zLP2uW
xoY1f0SiOhFDH3ADjUCIoe//N8VJWAL1mfZ2D5UqJ/yjb0Ad7tXvhPY16ZeGG4jg
p9PYnv7KVUMhV+1i1heoy/zO3ijvQpflvI7/gWqg9WlU3D3glMDOe82AVNfX9hME
d9coAnBRQZMP7hGTGmUc5dINA/VwnkzcQt1a7y7sDlppXVPbNcpmRDHqVQJaCRbi
1MD43MHPbKaCRMEQUk7qRk25/ZVi7GtkHxZfy3m9jhrLSIu9ByhXEyq2JVPf3re7
b5eQVlGFJaJFMcSn93HhVK91ca+JgBheXyQQJrsYpqwD7kEOnrE4jLmw2+JxEGsM
WO7iWl3DN69kQ2bZxI9QNUVmFubJlwEjR8LZ4bD1kL1i8RLsvsMA+UHVy81qSYhd
0/vzx5QwIgdlzEnPfK2DhgyFCRBl0IQQcNFq9IxRA42ZxJEhVbGonZqho3kSqXev
WmwfcsGvcQ6pl9sgX8dmWGpVkZhSjBlb3B+i1DulQ9nnLtw7rB/mQWqSlmPbXiUh
BS3RfmneS+fsWLNkHIaqyE2BAUkJDKfP4Jkw8zzhPDUn3NnaiFLo6yWn6I0k//Sb
kg9h4Piz/SQYNBsEYyU4970WDI78/1YvP6SIVDp4+gYb3PLirSeVuX12YLYllAFl
ZqLteQbxf1VVfQSzQC5tNq15d9XYFOnuDYrx1bcxcHLmM/n8gC7kES6tH9XX/FcS
zA2AJJwJ+FaoAH/JWoEvdMSUFuE4qJEK3HxF3t8NRnfakoDbWllUmJcjz17dG6Mz
WBIPS8PoUYNnu+4Qddm7ibV+wKkJpn3Uc36o4viO/5MJbc7rj9Eqt/QwoMb8qUDc
TPuTlXw6E5qcj+jy0XKSVcxSl7i6ggH8TVoozqfu2Tt0RnR0HUAFsqkUtzV1PiYG
Zjyft39ZORQO/AAG6UYCslyq9XxvbuxxwJxFE+1h2J4eYP5Q9vtlaWi4NAJpXlEh
BE3Q+7fpgcmSDpTq4FKtWbSK79zNfGYiVMJE71V7xrr/baLmmQPjuBTSV/hTi8e0
v13itgkqEuVvRON35kBFqytVYb8Ggv0z54gyx5ca+d/WtQSZ+e1+Jhx79xGJHcDQ
prChdPvDf+1bhZx5zfAqCMIEFPTCdOgCpXUrSQZUL+sKT9L1tj9tEuEGmDnDdJfW
FUgM0kJ3Gn5reJUBRLeaCuI2CLhoydR7+FITkfs+zEUot3S/0LsMb5eA61Ls0pOd
yQMuz6BrGrppOGrpI1LnDi4icCQxgNuRC+KFg24UGQqtYTcXMO+hy6xPPOoSVZkX
zAL2kUf+XoeiFayMYReFrmPOppAjQrJQgulu8ULLylyyCgj5Hw+6hYzS15klGTlT
Uw/8zOy31oKmuVuva5L6anoj0lUFE3sSGy93ho0Cj6sSkqZak5tKWbI4e76TyMxe
Uu3kCyHdJSggUgdqs/zL44/BfbvFWOLbo/pbLw7IvxHArCuj4RS3wioiHzlC4y38
nzG9svzk0Ncchcn2D6ZiFA5e7MGTPjPkOy2XaL5oE1FG5RFFnHmuQqbvyEx3oNMe
0lJpla2B1MXLOOuHIvea6ysFf4fGIPKV9DYQDuwPPT4VUcxLRigf8gV1d3lTD7Cu
DLryZAWK3ZDc1BOwG9VFISk4BInd3eUUF20C3G55kYm++wrmoSGhoRiTkEFVioDR
OM4qMvUeGlC5dJSbQ1VPs/tqoH3spghnXJXz6W6j2y4tEQ2fgrUOnYMcUwovF3MJ
qprx3feCQXdHTnSQFevL2qPFwO7LPAjIUth+HZVVci164Ahg7ZVAjrMEw7I+F4Fb
LDprxDSwfNqETk8+n/s9DLiuSgSTi2V9rVB9U8HUwduXSnibqK8NJkbdJRwaXX0p
2JdoU+HapnAaS8tYa8btTfNubnepgOWU8bCeorShLusYad/+VJkPuhn0KVymlIMM
1KBQUG+PEfzRWFxYu0L8UtndkWarKDgi+MvYL9fQZrbt4snLQg9XzDAeq7vewS4E
xosjMYs18qbJjDRXeXtmJHSULB2CgZFefx3FyWll9RVAzlYby8g0e+tSS3qKOIKu
Z+hbyFE4GLmHjlIyBT4q5bT7nzkIhx/amSn2oUv8hPzrTQMUbubB367mHNZVGZpj
HoGNvsiIWBcTwRgQHHTHgE3ytwjcdtcY1ytmQlVt4nwvTwdNuUSPUQx3KilvB7QR
Y2Sw1aPQeUKNn5uGGAB2BVfVtahtkQ9EnkluyvqKD0zo3z3nfb1/zy6Ws+9uTeNK
RTmyR/UadrD12xvtIQcshGLqnYZhtcPzkjsWl9s/naAnWgTTF+KzaM4JBD5zetBo
ZB1nOA/YoC1vpXdLQVOGom4Nklb7BHZ+Dnd3eGQeb7ubfMmOffdGRJiD0EkhwIma
OIAQ38eZFEREqcslgXkch2wYZWJxT5EWlFTJLVf3fyISeM07fpwmAzW5VsOg5Bbf
E+y1QXlc8f59tcJ34VPpASCg1XrsPDOH0jfn6kvcHgKKd7OdEZKxYJakqBm9mZSr
IHgeBbwfoSatDRJULEyptxsqx0khkTwa6JO39kWjTLP/dMFhM146Vx1j2ljnLwlY
L3nOGmySK4uPUGwY+Or3gGImjWD2C+MqFpYKbuwvD6iJRk5HddJo6laBUL4ytNE4
r75txW2vaZp4CiSRQgr1U8MrFLFLhSxkCpfjA6AzuSQBWRHLSZ5s0OSB62MpOwbc
5+gUulxifFSrEtAmlHjstflKE0fz9dAoy5iLGu9ONfhbNx878x6DTP++oZcw+OBS
r8OR9aIAL5oVkfvLAOyTst+udnd4Qf+OuP/ITrYaYEuUzPpCxcX+nO82a0tpNAza
B/OcVHA1sHJQqFo6oR8ylPz7SRVl13URmkG7+1CCR6e04diuw7MnwMLMRu1Fzok4
XIw6mdb6fQeEybxN3nxdd5QnMc4aJiG7v7szUxr1FamdkARBYc+2T8mZfS2zGhJZ
diaa5+ltspUUo2aPmhfFBWWRamASAd//hdC5sOPHfknfMo/NgR8SRjVDedJLZ046
8GegeX/lF3BsnZPy7tk7QMUlF1TNDEjckggXBwM+ZMBx07VK17rKompWKPJZxqlQ
dftGqsJi3TLHgdOhOu78nU5C13/+GGpFCfmYO7ruxU3Pi9c83cfl/1CmzVre6pVd
LEHjgRdQgqMiWGZU1c/G7sIndHgTkAUS3yzCU+r+tQHKhWXrC5Ar1kaNmPR9nxqf
CnhJ6qc0QHmBkA04xA1BV71GnedCLIIjP9KaI5BeRc9HWhR6G5vu0yWQuRb8Plj1
K81vwQMxvz/bWh6ijZktEeYz/P9aDcNFj82dKxGchCZkZYLDJwgE6Tc2lezL7nNJ
Dl2XNxH2dT91YNhTzo52n3AN2lBMqrlbRDj3Uf8gtCpu7K4hKk/0kK6SohTrOq3R
1AlKWo3QneIt5/W5QEdzOjdqNfd+fbd6uTCcEgiKSroNVtS43VHiBk1rotb6kXZR
cTm9r/DUCi9VITzeCvg0I4uivT2hqHsxEBo9Ppyy2mwoKZH2Jq5dcwJLDh6t+mYI
iMGJpwhqHS3uaorwJ728pzTaMIkSmtXwzkTKbwEDospp07VKWyBJont3N7semZz+
qKXLzyO6ZCw4IHcdtOvFDKLPCkrzvoThcB1Fc7F4d6rWpEPOW9fpVX+SOoD3HLcP
TBk7tzdL6xSuYy8a3uJex1B/52/BQHcBZeFY+mf+9L4dKpM7ManceJO/Ah1mU1i6
iSAvLaiGk3VgzV2eE1mp+RbFVxc1H8k9hbZmo8e9xLE1ppVd0AWSizBwkPP5Jdb5
aVK7wcaAP5f0rY622mzVO9LR/smVv0HHtoryHKbxUNUWRC5u3Vu/Jeh73hDsJWht
KGAbFxmiKrTrKGT5VEd+49TwtwL1RIW8zSBsLDQ4gkb1u1NMFHWtb4lk0erj6J8H
8kVxgPaofbAMkUP2hF71Ly0hsXmPb2fArrCmhrs9ZxLm+cTw45ayJ8fwJT6kgRS6
BbWYDPuBP/2ibQVVOKPIeRr/028wzLigk2UEufExUrgYlg1wmJ2MBg+z9SF9Ieri
dEjNl0LYq7FxileaOxPiUzEJqC2YgSwUAfNEYXEsoNNO86L342FmvKGvNBiynSHs
CAR9B9rMgIkLjwPtedfuXVovNEd1XliL74fqghjoAwdaWmLS+k+mrqCr0nY1dWff
ajVOxvSVP45KFEPGnsQHSQOe10sylbw2jv14ZNb65f/a7yAYMay4mn1jMl4X2icn
5515YQK5cOs9hlvzsxjHtB4DygsWfCjQSt+nKJTAuqVqru7RrIsKSXA4oRmnxyYE
wntTIxIRmsHvKUH8QZ1QPelgsgo7PFx0S9JgcBZzHf5ZLugC6hMLgM1rQpoZqwtt
B+jYkM7mHQ0PaAwjKNqiBiDcW4A5cIZfbjlm+ndmyR4ozxht6UVVcJBNf6UaC+ZB
Ipf4Y7L+nCVXj3c9bWtI2Dop53eJINv3Jg4+oJE4q2FKn4GhhJ46OeuwMTnWIvrr
Gn0yV4ALBi++mbhoyvxqNMLUjAmuGZx9pEe/E/k9qXesuyIfjcpw6cE3m0k2OapX
67nDf3tdwR4ko2pdXtaIz3HxUm14HY4JpNO8gjg/PUpVD/5cJBNIC0zy9bPRT1nY
iblBySzK0LDiMjTAY/vadHfQLpxlm/AVSAHIRSuiKGXAASCrEy4qr0i4RhSFjlbU
95o6voCko2wIZFt+Rf0xV9qHBxrrrQ10nr89CPh0LGsRsa5L6YAQMdkfU+Umj/i2
W7Ld6GllI3eBbHMdUTkjMSmJCUcy88Qr1XdnXoR//AWzRaVIU9/4puLm6t73lexe
UfriHCjzaOLue9RIzfUVhLWVOB4cZF9cTdcVNvfENSvZnhYZd9VZrOtIxp7q9YZ3
6rZj9w0+f+FEfilSrScy3WtggJVH/+8VhmnryowlaWkHi77PP+TG+ff6ROk9Asmc
tD9JPyiizJnrxohDMiPftskQVAEELRu7KYi8DB1ppC0RQ+gad6vMJk6rnb4lm7Th
yiK0PUljUlXH4qmRJs1cJgO9q0w6o61v/k20tXfnKDJqYIFs6aCGvqAbvTNWfaiR
bVRMCfd25cgJUVHaq3b313x2Xu5XghUW8CyovQzVXee3B5HYssXhkWg8cY032moO
S4b6kDKum+B6rrj/4J8eoGVVJWH7L2JGcOE4s1pJHiA1AQ5uMR65tmfSz4ZHV9ll
DK5fW3xfi3xg6+wScGX5w1kjaF6uqv6K7qK2DI7RPFLpsRXQe+03CatTM7J+5BrM
Hj7Z/cNkx1wvfLp+3+oeHTyq4N6D9KKkR5k/xec0NSaaZ9bxJGuDYkNn9TSia8ld
h0ouatxyo2Nfao6tlLzdBWgskF21QT3DES+RsTb7y0/Fs25c+TuNrBP/ZXEsoxjC
j4rnNo6zDGESm3Gnii7Ak88Hn0NkXHZUW8TRqBHDekcGn8DJjnEiUaHRtuwcWU9b
ikbWBfFJNt2GM3SD3YxGFFaFkzzeMvfn84yc9lnkGxpAKlR/MuU2+yYgDKu1vxxI
c4l6+jFmv2BkN7Y7vwWno/SnLuUglhy2AMLATtRRcb4jlFOndZSmkOJ84b2Xcfia
d5a1dZVCGBdwl4PcpRRL8tUDKELnIVyjehUeu7UzDnDV1fo2xgrQC+NM45RlDYmy
vThIcteb0jAmPKeiPy8PhJySjVwpQKXeGBx+ZwOQsacjZA4xbVtNgLpLj2V0pUy5
b/GesEgYqvfMoTRImzW1rm2VNYWfOtpHXpoF05pP9upxpXf3XGXM9SlYE6ML62c8
y5maU+/Wyvf0UHkWxoIm2dT06ZZAeOyQy32nYNMyBqs6EI7paD5XTrmik2f4k7HU
nkcgffmJ26df3wXpwmYZEZDSrGVC4ag7b4oPy4Sk2Gv2uhOzSzaO/gzEvfl8K/Je
0jHEU7ShDCPcuZlr5SE0aq0FXGTy6/lMSp76wLV9PBlLiljSmWPybSugob8XjtPy
xUTjmYnJLbx0xyyKh0F2p7uMdBmZtPXWnh2ah+OCg5IpVV4t1ZMgSybem4cUTs4+
mNlabNIjWMqJYGtKy5ZBpsYkdVvrgN63HLHTZ6ToBIgWev469o3lqfnC7SisvOdT
j+iumB/nhDDjnfkcS+cUj3nWQT23OXxr6JCfkcg/E1f0AnXJ2h1L2WBBGe62EP7X
qnuZ++sdEBFHklyAJfI5nSXFMeOcuCNwb40MnmgAthYdTjWASlEMjYSPqnlxYG6I
M7lNOGhB5GR1+8cJ0gLxcIJNs3Gj9Fnd7UJZSPki8UeldwK/SuQu3slPUDoahbSU
PAksSAB3oVjXUmU7yov83hBTgWOqKDp6l0m7Im0+cewpSF1pcFM25Fat1HBs8aYj
/zbIaseJMF5/PCtp4m602v8DYc1Bc8x5MBzGNWjVPNc4VfVAxH7/y4T8jic+Z16s
yqBdPC8UxEb2OdJneGd1CPcYQWPmf0eM0t1cFw93aat8jI6Ptprw/fO7iXKZnzmI
kb6TzxK6Ezd0ETRy8EuKjTWIjAKx+rWU8ONVVod7lxpoq1SMTrhMFIe0UsYMF4Jd
pzCyr5FrLcuRF5VQqapnqPQ/kQFgqPkiHNt5YSQDkEnZWCK+cXRUrWDlxRVFWgpl
kGw4HjDaHCWqqls02mbsDz52JFcJb8uYUEagUNsFksTBQGk+NTnn18IqJM5L9Z04
5uhxEkv5SMna1CqvDU5TWuYfJp8ZdYucmZuvpoIYjf8RHJzYAP9izu65B4yNAHtT
VpwJRfu9RMzRTepFp//0008JBo/XrwiQLL16TSU92y4frhYvNYl0GDyk2FiE2v4n
p1a11j7gLGQT+rvibRzWICMwHu/hJiujzCz0QWyG+/TS3xzgFZlb3fPePJkM6yef
2fg7TFhySaJkLsaf+pcHgB5/iyhRNMhrXrQZGDGDPdLlMaOc8w4GOvJMvMelhLNL
L4XhmJNRI9o4qPspUdB2D0/lX4XtEsZ3MVE0XmIKOTPNWaxTkWJEg8v18Hjly/dM
jy8GC5Fu31qfXOZyXQEOuAwhk+OI5SpZCSIRmaY0kSKCI1fhoi4iyKZ2PVj5jUHm
5jDH1cA0CQF39pdZ43Pk6wzuFZXNtUinOMTPMhF6fm8oAe5B5dT/YkHtQLB4b90D
Ss+PRtFsb3ibLbRi49GK8wxvasxhDsciHACXWKtMyq1KB+dYc4Ev5jYQ0xOlAEyu
Kf5FJyQxCwf+tTgdN40BLOVhd6mYUwg3CktgqT767Vm3cLOgswis6ecddd4019Bg
NwqIxJAybvz0cHhV8shEQq2UP5DOrSg19ZfFcXbmQK/Qs5/nC9mbTT9wa0pI+ojh
q0JsstMFE1zYoXlJSsIRY0VOId5W3uBtzR0IyKsqYmDy8jrnNP2ii7ohfzzdm4xf
g/5dr54h9S4S/XWA+Bk7eRlR+5kUdEiftZgKkykVQ241Csx/uRXhnvLqBEtmUaRG
p9/B0uSueNMq9k1g/yvIlAt4newEmyadite9Ma1rcO9lrf+xnyaG/SpwfVJc0tUa
Sa+TcFm1OWAIccnz+S8+48wBzczWdsQrxKc2/9Pviet7TD3T6xJ3N2q2u/O+HzrE
+oe1YkJOCIeYkcB26SriKPWe5S8GEhGT35xt+rSYyNiubIyKQ5ApUcqZSnoMXPBT
Iddr9t0klBGAz0yd0LePLOQ88rzRDo5YRAegQC0z/9FvUE37dAUo3TfOlFNo5OO1
QR+Qs3+n+RBpIMmL4VPSW8AOJNBL9xwYR3JMsqYQARFYKvPvsTz+5+8pevYsQYej
IqpQvroIpN+7McofVAsqR34cLcbwvuHQX+wqY3fylYFBuKugR32eZj3pmIvp1TNF
eEFozczRPUZHBxF2LQSVJ2d+7R2YApDTNRx2a7/vanY/z8K7pXnGjCxJ/vrFMeZL
sSbEnFflo+WVwsRRjiFdcbOw9K/B25YpSuNkMZ2206z1Ti0j0Ai/pDT6prMxUkaO
fVd1dCZBpL/srarUdGqVLjliiBmHzlzWr0Waxu7bCITuwmke/R4txIrm5tuKCyWm
JVG9B3SD9uwX82uBR1YuVIXWXM3C+tMpmbd5z4dwO1JwV5ltwJcACTr0UXFs7SeC
2qVCAaTvXxEoZvRKPpJLnxBYA4c1EyVc65hBnsoN2ZfdPT3p+ypEiuwNAyXmWH5w
grYWeQy0Fz6XfJ1J0t3366tvIe+f+b7WyHQuS5//i4H/w/0v4RI+RCgZD/FDlvIP
A3iLHh5KY/V+bpNXGDa+7/oVpuVT9gz48mhvnjJZ/zgE8lV23eJBF9PMSLMXYjcF
wP5LNj7gUHj0frGdMPhBJkmH0dkl9+kX1PMoXTu622YSh2wo7yIs9dxm+Vay3TL5
Gc16a3PPheZ9Vy7Zjkl7uMj+QhgyGI/HxfmfCOIgeexSZb7PpRiUtFzV1Mj5kqCU
Y2gh6jIv/SRYbFHNDhJdquPDWARn24JrDTrhHkbsAw0GXhsHUwKlJkP+wsTtdKWi
JRgcRpcH82SYMQHyfAv/kHRHbFAoUdpuIQ9RDHdaJJvigkRHu/2/VNHZ/n3MD3oy
ozG2rxwtTBNJY7pe1WRgpB3zPMXUKdd27uzf2iUGiPTPsvaB8Le5kZV8uX0fH0Yb
/SM7DPQ+JmBi/mEOaN5yDNrIn5fvxlfhhz5OKki4Dt7G6FC7nONk0VbNiEqEQFcE
A51abllXlsHBW89Ycu1HYOSBJEnw3Fau37cHiLab49UbaGPIT6Mw/1ZYtt1/FJok
2O6K3hjSShBxG77Me18KprbjLHDwlDZQ+ymrHq/s636nI4CzH7fsMHX8NvQGrz38
bEK16Z1aHBaUfIDV7D13pQSgjgff95/0zttxaEO1xzglJEsOHNCeKrXWmEHU7c42
hZN1A6m7VOegSvPNVQUKqhk3UVoUaCPNP4Yo+IRbLZE7CCz77HDr2TH1zfEnTIlU
bIAA8cIN0N8eKw9X6I8Y+1FzLTHalbRQa4lWh440nFAB0S2XSGY2QoITVJhdHQ72
Jio/pOVsC4RVBvVpgxOL+SPcbDTlAVhKYyURVhlbcnVIAVh/Rt6Bpz9srwiu2nW5
YK1ZLisJUJ7a5qwO2Jftn5la6jgPUS/ksoa2rgIpoEutQbvt8bWMkt9cFAVpfUCB
sFlemsQeeKDW7q5+qh1M/Jt+no2Pot7mAvg3DwCzyzMBXuz37ZvIUBS66EWvF9J4
eo0Uk9j0zef/16VqiRJ2w6JSC8m/EY8yhhO9biw/UTPh8fdvSM1L6VR25+KYzIQM
nKWcBjbYKL0NVeup9pCPRn7XCJLydOF2x4dwnez9QaUZnuhCMB3LXVGloA2mqD9j
NedcgWV35XbWrK4zjVOpKWhtA+Jdxf3eGGe0BFg4AhsZeI6ztcPvmu1YAf9CNNtP
RRLGsZwm1rtlvVXnKfvrbt4CmRcl/zFoBb4GLPfYzsNI02V7VtMj+gfYfBzpFKcb
GWoFzGFZZIX/cd44HrBaiXIjT4t1s5Xh/fKDJe4dgb4wpwSOVwI8SlQGvT0bboeo
DuZhHJLBcBAoISxF+c71Cm/gjLdnsszMwkBCY1e9HHjqqJGZCcVOXG+Fq3uRFZ7a
r4lY8De4CSDEWneQiXOmgUAt4EWNwRqAQm+UdlZBAocqWOhcKVNfzuDEEIww54+G
FSe5GUQxeRLo0/M0If9PxEDrD1ZUYLVYJXHMFe44cJdjlqySnTqkDaQslQgJKIeF
K7IPxF/OChj8zG8slYdpxsM2jp10viH52IUqnZV8Gdr/B6g1R94EsBTvqafl/jCY
/AbwzxeEMElkTYMzntBYUA3P/MFy0iXh6TIF16yXAzDtlxuKshRsiPkrOo3AdEyu
TPOUp4y/cNFCLcaaiIEEb4j1mZC9ntvJL35E4vxYAepIODBKa+nKcVml0xkmQws0
nrxiJgrBkGKxEaYFnqfqqwVkG3V47O+CGGyJCWa6w5O4N2dxhlKtTB+tSBCMIo9e
CnXmbv3C9IarF8MlqB7MQMKQeKWndzYjnFmj/svDTpeJ8R7hi7GxX9L+j1rqthI2
Cmy2G5OztMapt2IdRYwmupCVf0asLnLtHL2Tvm5RGEGLRosYrAGpfRDnlbzHzVcJ
rmoI+DQmiJpxYZ7/KSi1jwDVkJ6vJHFWX+AjUL4FxeYrwAfkMmoTikmxSBRGSdSP
el76gj8ntbkaJxbxIAZUMG42pvDayVaqs0DSOZx9Sa1UDg7wcNL5MldAUXhQcksB
dh5nwe02VLmkOCzYJu7LHfWOymfw7+D0s1fD3p0KVZ5Z1j7JNYNLGzBf5X2xnNJY
0+y453w+34kJvBgNxW8Nn3XiXIPvDRuyntIovV2gWyX2vg9fFS5vtHLSAYwg8Ytd
F30OkUNQR6BWozKzjHrevZ6mX9teFGrvdSopvFm6hZhhIeO/Ts+p8ieh+hxYgWXb
QL7uSdiYIJj+GV0emMyNqjNqVI5Xe9GkpFXDoub3anhOocQazRYMGOLsYqtktOiA
9J/ZQuMgRFtrqKdhJI4EmjxfmQA2Fi/1Mac5l+eJuWyCD8zRH+IUE67NSpZlbGbR
3Vibi1ZwXQHO+/jy5OJM5PymE3HZQVeaRZ63PIVisLOcemC9ryuDbdyUkf0PlCcD
vFJ6Mw36DUzdcY7GzGwoJyfe69CfN4xHLfc4ZFUflthnstGZLIJvfktwoDYGF21h
5HSRjo/B9Vv2bMrrpptn10Gtqoeqoen9UKhOSVgS/SMsD+doWiQkzewBdwIMxCIX
vFSSlfXAC3YJR0zH/PxY9+Kxxbu9Ggrk6TXYyHeEdzWxIH0NKOB3FC504ruDNf41
OOlJLWJ+sEwEWu74OzPTpDUsGAhynGCkGCXNL8GxXvl1Lwa7gKR34UAu+ggYmah2
mtT4A8fM7aIlCz3aZNFJWC8OjriuelU46pnYNmiIMBeCYiS79PMJYsItfziikjMx
TIpjenGBry05JV7lWCVkyXWUN94V1C2imZWRhcOTUwCqec7+VXu/5xoVpZTIETSd
6ZLc4fON8SK0qnQOZ4itMUScWKnru6QiCoCECNODsAMdMkgFIFTjVuCBHZCoElrN
eG5mElTo6/DDBDG/JHjpclz7x7fiVyTTESC9cWuyHAfl0D6ftWT2b9yAsOal9oDk
/l0Yra8/AsKxckiaRSjeRr1O6Yv2mLKXRem17idQkWzP9wm2w5bBzPkggLYSiQgH
6znSnsorJDYk7uzNdfr2AxOOqxG8dsDeINBvhOPeVjOyvBrezFy2CjPLSLLkJUfX
1ufQhcQmcRBy//fTi7N125aq79FH6Vl8Vs1LhzajceDrT50I0pDFkVt4Jx0Bjifv
LhdaS5SCGPzqAANpH52V0q41K6n6cQEEN0goNngQafcvF6vS5pos0Xje553iX3nq
L798LFxk23ri1E5TYrj5VgZQ0yUpEhLUWyAdQEMb31JRlHsRlWyQvOw0YmFmYVaP
H2S/Do5MYR8SpPYYP1C3R9DydtNFer1O9LAjfs5YJmPbbBJ0STqbqg7YMTcpar6q
4jFShS9rauRepcyKhJcDS/gQ1JQAntdTJVRbNy4hWWWQI+CxX+kd6mAx9jOV25n9
wW+ydqiPI5QziFp0TZ+PDL0KNHw02s1HeEsoUq4eZe7p9nm8ENGbP0xsbm8FIBqk
/fqMXTnD1fxuPUAHeHzctC/uTdHnjcSOKdeh2MhvfNlzFrGf3xTl5J0MBmACot4L
bus8HG0ueUBDraAM1O3Rs8NrZ16ds4ZtlwGUr3DOeKL1OQg3rzynleGLVFhH49i6
jbF7Gf/ApBQg4oW77/078LfjwU0xqByvbPGxNZlFT6W3d+l7JA/JKzuO/a/vD3Zi
Shy4YxGi0nrSbriKjAHYq7m+XsswwYGq+VxGO26z/AAreEDBZDhjwg8lXHSCC49K
YwQi1Laons+mZkHk0mbT5o/SGy+oB11s6ZvnpY0Ld6Lm0rJz79vWOm14wOdDI9YM
2heaovWuLp3qHE0F671dqobOoXvwN0d/hCp6fhN3xZ7AM7vz+7/HKJkiuniLlkw5
AZm/IcKFuEEBVNeNr5qkazd5ByReLwyPfncErfuakg5xOtoJN5+rETQzoCtb6xo5
xP93ABL9Oma2P7kCH53+3MeaGdGo5bxcCL/I+SNjp6npo0gfE8UoC6dp+IgjfSH4
83hQqJKrqNRVjxdjPuMBHeyCFXOR8OG9CWzuC4KltEKRkTQqvRG3hHfud5B0pwWU
hcW1p1epne+8GMPvKUoV/eRN7S8fENQsqpyHuubzI3pbgR8qOzJnEZFGlCwkNiBs
ucgKLWE0W8YCPI6vWSyhdLaQU3egYSFaL43cqELojaAI0B+KeKPiP/K68d0AjrsZ
mflgIfxnsQ28cPKAZJzj7U/otWLuOoD2CK6h6z9lfZjYzSkJJPG9TNNtC/6Uabvl
VNfCVWWCNiP7hlid6d7zX6WJ8aHWltwTvkK6PHNaW/vcmouGyboEfkArbZHzdG9c
nlgbtAnZYVWkcE+p+ztV2D3EIYdK+zqujDkk5RFaME4R4ncyfeDzTfJaBQSyp9WI
8QE4DQ/Q6vPllNUrXi8IuxzsVMEhL80H+9vs5q1PJdYgGBI6w30pquRR/c6fROFm
GKLqF/hV4PXphnCkpR72i/97qc4mNw/YrjK2GP5/1UHVhYX/22HdJK19YSVVFxmn
rp+FIQ6P0ufzKRRWnSCgO/LRlIDvGTBEoJwaqnuOp6PO+QScVNQ6QBEcS2n+gwGd
oNOjvTNX2ughj4tckPT+bD9CQhWVve7EldNteumNtO+jOBffS2WP3MzAaODiGdb8
6Gsgd4IzmD4a19GpS/2Y+lTBuB4OBn7U0zRNKMQSebqlzmWvbXCMvwyGJj4c8won
/y5M/Izwdpk7I8yvkrAltIjglNbxr1V6JNFee0TjmSxc9+QSKyrEsmEixKEjZ1dV
+i2DMJru0ikwhembnFMepE/HEqwS5JRS8JzgsfWS7SBoIZAiU6rUpWblRqpbR8t/
sVTAN65Lm8D+dZFsdzV2rwRkNLiwPqG6WyP3T35F8ANC1A3gK69m9lfpCV+uW/e6
3AfK0lJvmzH4K5mpTqtL9Qyd/el0EL5+jATm56kNP+B2cEmdx6Xj6YzM7oDdJmbW
Gs5rCOZYZC8TunMU6ETUCu304XNoMiABymQsQEWJPq+p7LA4tRMgClvSMeFC6N7i
77i6l2WNswjqqbaKV3JyWsegIcOJFukR1UKB9I2SW8m8DV59W9jSjrLGR7bOQRM0
J6JkCFErwZfa08QdI9q5MetLpKiqL7j+tQye7Xqz88fnalaQ6ydVv1LrBGRYd6FC
4xiU33VDKg6MYN4WtIGGc7uVXvWXvzLzz8SMxdPNLifR5HGBDQMKlZ8kecXZhV7P
2/m0UOaF5ZCmU+f0cLo3zGE9avlrIkVnwqjYRwzxdVAjirn1GPiluVDUe9lXE5Sn
8hzeHrPJQnpnFLdKMJpPf9DvJZrFqIJaS/Q6Mhegb+u4ZNmLjbYRBFR905pG7ggz
A73p6I8bMp0eofbSN3Z95wzoa4rhvPFBGbog7P7x3oZr6YEwLfGiOQKA82OnHkIi
FX2OVB2dbe8rQ+5BoCJVnfDMR5kAUps6Ym8noP/gyyYiuZB0eBuWDK0OHxLtKpAf
V6oC1q7svusW/Pe/0G5Os8AWPNdB+hRHIzWHFMmxPJBfQ34qIBinWjZ4Er9eCFdU
LZeY+AKrnv4Wsq35DLMIWdhOlS6om50liRRoyjzC25CSf+LZ40iUCnoumWBkV17x
fhlb0ughy8Ul0g/fnfS0iijnmlkAWHBNhjzc85afa2H4RwWep6KAigSeX/HcV9IK
piEDZbWZII01bUjn4M5tMs5Mu3jRiUTzVZKY6ZMHzJIIzl9ze6cyiGyqIkPSlzUF
IGkZp/isi2liZb71mSZ4VfGRXUAb7gSbaxJ3rE66iURzjix/xDCvid7J7I1qFoBh
vhM6jOXZY+MfyTN9yChjBYneOA8PCm5lMyfzSpUIsdJon+/O19URgrPyaOpIj1SC
nOkeaY/jLeyGVSfyrJgR0Nt61o7nsE8UYPKuh4ctP9dS7OTfrNcM17JblHW+BKcI
ZAoxFyl8k+s8TAEocgzM2fWFm+tTizD7nVFcUqVjTOA9ud/d9fYS8KKRplNtI3NQ
+6yjy5vcB+3axKwgduuYBK1YMoPlenZl1PbVaNIi6FqzZAWdTgj4mcsXVd4oxh6/
perOyAy5o5DuviDnt2kcITusa2urbTyX604gkVNAwWfUvDB3KuaqK/t9cPLXh/WG
UmFrN5o4rONvVc6mqho8IApkhAzoYxIuFSogyW6iD9LTcuIEXEGcdPCg2vnPHslN
FWyvYd4v72JEAdn63Ayb16NV+ypfnU+5NW1KeWm6aJtkFHAcbzj/wXM/u8hr0DD2
EZk0sd4y+3OnLBQxuaGpcql9aS3Dd9M+PMqavV/gnYStkwAEI4suR6EVBf7X+wpK
o+FglGVhdZPSSioYzOrPFSOhyTeB14OyBi3xJOCdi71EA/u8Ob2tYUMy0BXUR7zI
ikK8WE9nB7orPiZEZKzrNS5xzBgEm35ENYUw5MZDdGOHQBWaUm8EwarL58orOSQT
G/vVPQccRgvpe9S8Ag+p826XG2q6XeOar6CABtY4gS71wxooT3AcBT5XoMEOe7pu
DgZdoYt46f4TLVBlWDnblK1ZFSQo8JDrp4aBAbwMVpXrGYV12j6LzvgnScHu7eP4
OqCeWov2UbW9PwSRotcI4DfvI7gITNnV71hXgDf575vSHzheobHeq1nEFhcPfPoU
fk4KXXg7x67m70DrGFmbyPc56I3hEBW1D+zmMGzJiBRWVqQlsZ7UcEM5VrbYO0M0
V6Pgm5e+ObaYgLztWD8gCT7cOnmMR1uUy8pIsIrAipfEhIM+yzSuac8C5tIeVQSc
ecXWiP8IkOpafitmYyHmT8CA8OEfSjdc2PZ1Xr3+P9WyBMTvqP/zNOLI3+2KMJZ6
YsUamZ4f060dx/Vc63baF/9nWgC3UyYbbwxCa9L20qs+WYTr1+ZlPfy2OfUvxSos
axAzMuMyb32lSTNnRDbM+XqOknG5hcrTul7zzLPuutFLpt1t2wbHuQGxGYs/Bx6T
C3OJ7Z/X4ElYyR+qtRB+mB0+QINW5b61USGk4wxEQKpU83bDp3mgI6QB2tg9UGJV
JeMGtlqkdHv4gW8GYGUf1IyxrlBYBDjnJ1UceVPVsrzO7yPUsGN8XfkfUgJyEtat
u4EO8MZx0RpUP/y6sMkS4s8n5wT+elsynChc7bEhRO+uxKGYIkd5Ww1QE5QaPfo6
43aF3C316BTKnOZO/bgEKO1DPRzIOvgG7J+s2afgMMoUscV2iZ2U2P24+V+X0F3v
jsHQrQeVKZa9ysb9/RwDhRyRpf8iFwj35UFH8W/Uf3GtLe8mTvqUcpIZ7i11Rqcr
DfWtAPy7w+zx3XQ4IJq9PK10ZSo3IaX/giDkx3X5BgWP/Co4I7WkwOvtLY5fpgdq
31i4BNOEe2OEJxpz54MdpzQYAyrXpSxDrGYeA6TAuaLbD7nRUIZ5S+p48Tk9i5+c
oQYxCrfQ9sqJfNE388/NgZ7JPWf/5FN9x1nj52dwcraEa+GQg7BL5ebh+SaSvxPN
LywxKtnbf5WPTNKvVIEL+a1dk2CsIkeplZ+6Yuqdq/mK00nZZ9YoBDGkN2U9Qlt8
rzf3SPFBbAJ+z+ImExsIVd0e+lQ4ejHc4vkyuZy7qyM5kB/e3WdtRqIrvl+wkfsO
ixwX6Jj+93t8ayYcNIPu+i3oDJ3yuiIAMYNX6WjmLf3JBNlTXIUILI4ZBBbnR7RA
yauWUVXPLVCoBqYkxEvIdC03uNwn1HjwVhDgx55CsFQ1aTMETDZHgLaY5NBtTy66
xfPQr8s7SfTz5jfIZWCg6XD641x6cQVxKTqTB8tXb0xuYGWruqNiTDyHy+NwxaBS
uqUNMN95agPNZ9fUbwU/cmSHQ11dgQtm+MKDbyqT7wTBAw9jLXDbFnBRIgbw3Gef
aOMAugU1/QQ01ulXkp2W+87Wqa84ZddKs2oBaGWhYreMgHJLq9yM8SokH+AXG6/q
BjRZcO6d/6CLrY3risRKRqaLG5mB+iRY2ulR1AFM2T8CzRmREmpdLvRJydj2kf4/
klxhK0rcOcE6jdpMIl4T7aW6nkfge83lXjsKe7e4i3Djupwr+mpW7olB+ERtf597
ORqVyuI6laXp3L6Al4xf7JJNW0Cd2WAh36Z4+q2feVBX1sEKdHwl5g83q/Bs4cpV
Lop+0VreXKtHqkIjYfb9+P6+d2/Dpy2RnA1TxYhh9ZPSgFr0ChYq4E9E+7W0nFzQ
Iaf4gfBlpm3Ph7L1tL3nfrttRtQLKkJPsfM8ABIhWRmoGb+t3A4NbKYvD5I+OXt5
DSqfka0BuZm85AC5Ts5cm7Hb5SqwUCjRO1q3UnyaqfCXJux1SZNqOYHy0pVHH81N
CaCqyj7QV3bP+yS7UUm+mgTlpRW1+g9/QuMGsj+VUGrWeCKDgFKNDTeRP9YaGADx
38RLoWiauF+K0w3EVxu+F2gIVWdO6g6S+gghVf8MwnEm6B6jE/WIstldomWrQogL
pfjqzudaa8wTJX/4WnyFHgR1BWk7ovn31qYbcvpgS3FTFE9KDgUAH+KKr+R/Ogfw
RuDetM3MKyzqAfGYMYB6h7Fb6sykiLcfNxbpnSoivTbNUVMb97tqH8kR2IObIPK8
EkAj/sB/zqE9DWG+L6xHrNNn0SRfLOg7SYY0Amce9hbKslD5IK6xoC1VfWij4IL5
SxZtuiX8+mdX2Jo4ZlKCzNI8Nxs7lqA+o/2CSkeWaRyFRazA2ljCwoDkocAmOwlO
cn2uOqfW+k4ACsn6EJL4Lf+ZKQyp2VXKT5JPbqMa0nFRYnnGrJOCJcjo16XA8Xgm
FkmA/ybARxJ+z1X3BeMhe3pi1t4DXYPxmvOJSkdxIkZ6yc3o4k0xwLWUljbf++eG
dyjwZ9i8kLVlrEhW9sfrwtDJF3AcYZu8pBftu/lbW3MTjQKLFcCNrWiPi4eiuDTv
p8qmALZ3+Ly8lvk6Xt6OMrEj9HuV0x/nVjl7KgAnFEMjsatRWuT7vReLCOP0gvA1
j0Edc8xTwa9S7OOssVt0eI99K7gOK9Acp2j/wICDOGNQG/Kg9Q12YyN7WDSj34DB
ff71fGKQalrZFsIheG2QB6JkMPCwLEgV8vn6Wt9eUBLFzcP2XcXYw1JUbZv318zK
r2+yEQNAuD0KvzutmWnjxDXRhnNcY0N6ILX+kv95FCCFdpocjyYS0Zy8KzXkMwsY
iJxQAhq8yFSvQXad9Kqpl9r5SLmETZR40/VgzeasTjyTv8EmbYR52h+LzI4e4wCN
jj1jJXwIzvR9vy+1cQYXQGFwCl7ML6bNC5xA1A77cANha38W/UDagCGcbUUohSg/
7Mpub6tXjpfydJN7ueof+1dUjgpIdQCYtLFjCeHnS6Z3pDKrYpjVJgCc6R2AVoa2
UZI1X1V5G4fGXiaUgpaf3JkwaxUooIpxh2GR33asC8cQYmDq5t0zbaLIqnYrUw3c
K9lN3maixwrsRrKKY/Andl6UP9GXrlxvjt6jwjxO+PktAuqC4WHm/WGLVTQfL9iV
CSGbwXFfwlAPbaAVj5pRzAKKEEtzEB+YTxLfX45rj7bPYt/BeVyJHxXvf8JbrW0b
X74XlLZ5owlijGl+nCl+Jbt3hujFaq+XwzHgVHyxlyLyLsQWxAragcWN2x2uDuE2
+FAe86LG4NTIvrP3bycnkvaOvURZCrjjgNZnnTDRbFksRGGysIBqhmNnfKs88C8t
lJ6UkWsjs5YCjrosgAui8ZTGXHWhHQ7HEgmuTArNsUl2Y0LR5uhOQW4NreaIj/4o
kTkMLPyGNeoDKGJF2wqEyuvCGtnu2o3QZA6imfdF+2ZzAzjbzRknd0+3L7fpIWd6
IO6H7dLQintQ9W5GxGePGc9TgYY8LUDm1Do8iNL9xWNMePAp1Ui+Fl2p7+FJ6dc9
PafoEqc6jF2s/LP7qgg2wvrUbX3VFW8Q8X/M5pzpbDgBBmPVeEigm4nMr6ghIm7u
jR9Z2wAOaH31rSq6FgrZZ0JDuDj8IJOhBfN1jbdlshC8mMicUK9lM5V4kJIKjA11
kcKDnARuBXbX8fW2cfliu1RvnO0DYesG2G5B+Ve91Jv9ZFjGpBj1jqaAfyNNKO5n
74h6SFj1GtAeY6vxx/oYkVZBFeqWRs6vLj9S9EubEYI/Gkc37USRlSAeqaWgc2Ym
Ln+LqXrYmmkj1XLe5vb700xw2aFVJNay+z5LJ2l0nCSxaeGsJMg9jv0UiBIfWExJ
iKtkV3/Afb5xVUbOs741661CGsRP46T/zxZTgtyQ+/Tylh3YqgHwOplHdkoyPjMs
yKpaSW0bADPVvRxkLOZ06rSvU269GdbevfWMXKGq7+rs8UGQfM0ddinEZUB91yzT
UjzWht4l15VIZXJV3KCq4m8EAjihViEnd8ofPE/AThAUPMU65/G5ffg20xxR2Axs
aiATlE/mN7bIRHAQ7FIKKOZWjYkZWIUlLLyDV1w6d0/bm7/6sa4Ln4NP+5JqkaJK
8no1+ALQkQKt3GfKuHMADefjcgq359ZHIW5c26pwS/dA91ZI24DmCl9FU97iUSwB
s7fO5SrTgfhbrA+44m+xpk83KdbRE5DAzxxMTvxzdJPh1+ega1y5xd2vSGQVxJja
oOfkS+lPh8G0McB4o0e0eP0ufMnpK0du52KwZP/wBmH1EbbbFKXkAw/0M+kbhguD
hY3H+2ZlWWRyUPMGuZvdaJosh9nS7Nn3FesGglqN1uqA0TfOrcmMYognSb49pklW
Rdd0l5jXwhE4JwfVBw2gu3Yy3IPamXnQ9kRL6IaMV8xz4sU9l+4o7ZLnT8y547QF
J3gQwoEB29y23/v+UNgJW0it0rxSTILSJiZ+aDydRswVKwFVHw/nnUJlD6XXRN8p
XfnflN9yt+dzGtLJQN49mheTMC03WgnUj7fEbJpGHSo9OgxSI35DfqUP7p8lChNP
O0AH2wizIWUDuiGf7wuAgq7lXcbmOhjynwKS9w7bgjROF/YbZOsYSHx4dNaW97DV
ukOx72BklSodZSVXhbdsK1FJj3sPAyZs/zIUDM/H/K9YZGqlxbAV1cmrqo4WzOB+
WTPsBgJyqzPXvupUhTxNLk8UE62Nahz+Z9yTGdF38ByOazeqqNwAZ9qiEoTPnNCc
MXaCGXU6AmcI3N3qkpqd8sdh7dyMMDWv3NbQMIIZtsXCGTeIMGDEvorxi3fYfDsP
DLhD6vFcbBriidwhZ4b9Gof8+Pg12liljeBKVcAC5yosf5UtvKgHFnV14cP23LrE
aOBu7CjvaReuiWkc40hGPVnK+WVh+GslS+CPW56lrwsXBQJ0FY4Mce/YI7XlIp5h
er6B2IAQWLCC2XDtHeuMeGaGactVquOb6nGPFy/9uzKzZ6fqOxpJAWK4C418rvk2
dod/weShQJTMu0R+TMij2pjkalgCOl7kalmhOFojQrYRL+QgbpRklluUSkfFTjap
0726IIyJ1ixcpvJ+fOng+mvLLO6Bra4kfiVnSTJ5nZ2kA30FAsCthUIxsw5vHMCi
9LOVf3Vz88ijP8HqnrfWZvxDevEy7+tfe6MrBU0HY63r5aoILFw2KPq9GUrTBnZ4
QudoOwNGWd8aK+ikUX5++XYO3/xEzMEfsKTKEU7q0Ufu9HMWN6dUVlGtu3g30w7C
IrB7vz7jecb8iEUX9YLj3AoQG0CYmA4JwNRTMFg/rTCtri/v6Vi6PuQxnnVYn1En
4rT4YdTy/70st202SXHeKzH9Ixi9vL7TjPU98uiUkBf3730G8AsLjXoc8HTyvtFl
CnNIvRJ4xkVXLIMqL1jPJWLB8bKCHJFgbCEvRRoSLM0acVfRcK71wQ49TI2LUN8G
WbFXLR6okrI7I6Tjl/t2BF7b7HXM4K2Fr5uUZbwSbLFkZwW8+gQQksxc56tiyQnm
0QzEeOx//esspuPUHq3+rqGNi1v/PoCLxTz/wb2WmGsLv78oRlckzSfmcXM8doQH
tLI/aMXbei4PwK1wBRYQzrEuwj/DeEJSPeUKoaGZK9cLwvFUNktpdJ+tQbb9m1fr
hHswu7E8evuIroi/sMkaeyap5cRnmjTtvUIKjQGnTQdIVw0Z2gT2N5Vz/H9F/41D
7vyuxsibq0CBmh5Mixn3CJIgSz2yimIXaL5v/Bgmkw0fQ6NCUoNOiS6icsFHh4Ui
vO6LxJ+re1m5y5sbDBAmct2HuB0CAbxVjp6reEb2gEDWwMGN3L25MqpOox5CqOpX
OvNi/XXufDyyPaDvZLd2boOIW3jiJQvUZNALOp9QF+NHjdzRojmP5pEhdbboRnvf
fe98VvW6/rCaUX79sLrnzD/lAu9jnMgR0OSJw3HWefe7ntBnoXAugbXJZI+cFK1P
yKZ0m9iGS+NQ/Q9NyAwdbLu5RnMev0RWJVigAUALir5lEPIuLe2lsDMG484Hk6UE
OnM7aNUJ5e17u0jsXTnw3DV3Yc/s2F3yiZOZU70syuZDLiKK/G1TQpcV9FHiv8pB
Mkmx7todiYtc9TUJIMj2AMk0kLPNxVz2yijKPyEgS9aorhwfi5YRZbWYsNmb7RKu
uQSPvMwuSGS9xpofPeYX6liTJprfgGylnBohESopMV2C2Tgby3vfJs6QdZar0qZV
480dnJqEGonV/ZImuadZZw5vf8ZQI+fC1tIzPgevD/UgUNxktIAyVZzpEbfURooo
cjMJJmokv93xJQujMOdosrPY5GKMHQ99wLVxMWhfbuVaBhrNgdeNRLgHKYFMu9oU
RDyFLBMcxebkCf+xnPKPfGahi+VPL5flvJkSRL5ABWOkwBq/QTi7CcH3IXER2iUk
2tZ+g4qizC3tpNrL2GgqzZeMTUOB3ip+YSDTQfNmK1sT1pgb0NwkyrUCCkIDlRRk
7UV5t/Ongr+tWKkHYkXaySCl4O0VJJKtmjkozmrviotP/K6eBjCN5EnPi2YVMAQq
Roq0ivLgQ7EYMwOVOCxxOUkO9bPwn+z0zeKlyAZ96oVUQYOIWvC37bedU+08UTdU
UlED1g7Jk4dbMfey4BSzB6qj05Ur7/RwNjCjy1/Wj4eD0pEsZIZftWMKqa97PAVb
EC7Du2AfXy1ldlfICPGXbAxe+qmthCxB1yJYakD+HpeZTb1EuwTYD/n5+UKg/Eim
/zkenyRlYF/Bw5rfsBjU0P7ewcI39RKJcd48J0UzQVjd4kSgMaYMPnbP8o9rFZjX
1ZsYUqylDIXTnPLYPOQ0B6kH9wQcTYA4LIrDzMr3XBqZQVDslnYlzqesVGDzgWO+
7CAARrN/xIppuLgAMmK5lDOKyRWJr8wk8j28WBhn3tOZlwAaYT6f6HRVS5PAd+zt
P0bpyZ/9p+A9sEY2CEu+dNtx5I+MoLadoUDwPREb0ZLBt5jDr3AvQ8DN3n1uqpAa
XVaPNhm+7+zwYIhaXexzQbqPFKYLlqCSDWyXa/E1Fn32FTuQy4bvvef4RndmYE9M
qxEFLkL364pLVH+ay0qpsAN54f919Yt9Rjjtr4Ps0YKda7aP9ieGtCYz1/uBKSf5
H+lid+Zfz0MJ5yVVuIxXwK/XFJrUwGX+COElek+CPKyWYJYazLxmFbXuQpHwTfSW
2sVm8wrHDoqh/KHFaOEBABQ/2oTRZVe7EwKErVachDBb3zQI+spB7jPm2Ff29HWE
wUllqRRZVorBY2ZsKFaMXfkXZ/Bn4g9YVMW/c9U/E07wCCyed2fxthi7+G7sTJ64
w0IR/KnUm//a+xjl7lh+rHF7hWDZvAkm6eq8611Y6mEIL6ZVwUTLKmWUnFHAQLLN
Yg6cZd7w44kwLRh/MrdVMFlgdC2GFT665T++eM5UhTl1aH34FyOPFhUmu9jfQExU
6S/TT63kw+ZOu2gCw6oi4Mnqtq1CrwGnVmmhM5z717H6o+eeRkH2nh2q1dWnbGDD
xTA+cQLr+wecT/3TvwKTjOBHn0SETQZKzGJMyCt9SP4AMD7nNRJtUyJY9SkmAkNH
5cB/W3HgxfKRuqFokJot2DqjjBWDlJHEQv01SgxZycCfsTO08oHz8flk+JMqmaMN
22i5btVxpj1giqUD+MTIjvZWpb7RREMN54y26ErnQXoSSle2jCgHYPpoBeJX6pVj
WMUXFPWwHGTGuMvHN/TQ8AsBmtn1YDj2SB9I6aYarJoWw3XJq/NOS6MZ+WROgWs3
BIp3X0+MBcHVnvbaWvUJ0Hb86E4oarlTUnSf2FELdOeUIEJNhctIRK5tZf5UVARC
2l/RCRblw6D+jPYABJSq6TWoQib+21JlBD53CO47hTm5p/nOcT0L67K6VVaDq9hC
5VQ2Y3NcJKboWMZawDXcoWbVCNAzGOEP61yXGEf/7fgdOQFmzJdsAEXHyA19HUTm
P16jzV2JhE+tvEN2XD6VcuUp5OymPFsxs1sB/thZvzUSj+k6864ZxVf6uShK+XSr
dsvYTFhS8jiLXsL794aqparvyJ8nL00fyFep2zYAPTNUqbeViL2flMeNcMsli1Q1
2E5vICRKuQoNlNv+qoSdG1OBvFypzhDzbA3I3u894BdhsZr5WiQ9eqWFBUrV7XW5
VBVo9vqjF72FcIihMjSkOgKnvdEhDNxtwbBUxvZvFUbd1XC4AUnMMJ+TcH8941ma
pWHLL1njZS2ABBRCPC4/tcXBQvkboSEXfyCpGx2hInmOHwhYe1mBR6K2r2nKn62+
jR5vJCyw6PbNaItJyFCSSJb9dowOz4Rqr/u81CHtPMut2xZcaWxuiixor80Gy57Z
KXjBHIWHFyIG1brS4CoF2lS/5dAMR4ItO5dwaoxgMcHiVjko8cgd7CUxIo9QN942
dI2Ba3wUz9PM/JGRnDBrRhGYUq6jpJszfoAkqxPgTpzKivjgsCwCfyD4K4zyj8nJ
0BmP9+8KOttHP5/Ou/shsRJTOXLVQP7Ni6pYalGXKGqaZlLVIO8rHDNhNXFPcndR
t9b6a8YbEhKEcfn2EJAgdDu88OhPTSKjs1bLkS5WIxQ9gFCyPHgAXMC9tngkL1Ye
oDWEGTyt8lgpG58sz5kS0iVDtQplfR/btbu9J9BzXALe1NeDejZRi4EdwnwMvkAA
LqcjkeFwA4QT0rb7PxX7boUrlRd95Nz8kup8VjgiO1YDEJREWldbnH5D7BT82rR3
usdgNvjL18rC3SR3AZfeecgZvMEEhMTpDb1b61IAKb6vLeMcfUSLjKqr0snN+79j
K4GL37mZX6bAku+touWLBO/az2zzAO2FtslgHECrG9oi/HFDrt8qCEe40+wx+tG2
oqbxoeIUjALyHunwr5ANxCpTbjzSjPwRC4XHwdBDIdj/V2Lcm6DWpH6yFXq5qS5w
jZ83eJKE6XHBD6ALNb/FYbr+HWSKfscyjhqvIBrqlAvFwRsIccI2JnfoeOq5COO7
cg3vSc/rXJUk4nqiLUXydRTfEFGzxcmZV8PWJrEr5t4/kp9F+yrr59kt8GxFgVds
Pac5ABzaoUFTEJEKlEiCTkeQCdoJeeXBmeqEA/34rawZVaCpCkrL97oHcqXwgvE6
cNKlG6DM1lDWBX9OH5Xnj0VNKjhJlnNfeLeMODWDY5ncg1njseXci//X7O1p+0is
lXVRcZs9fJ0kuVKS/q3oepRKk5F2V3fzen3WwTBMMKCylMOaAWHV2vEzHx4VlD+n
2+M1V6AiN0RvxEssVt0uFsZsHSQrJjHo05NJz5BeotnixmCJMxtMF0N3oT0saLro
68uXY6e2j+KexT3woW5Bl+vEAjvQ00TH6+r2WH9bXzgURJPtdNUieJfWFE03ULYA
+YwHXDxIDlqteQVL/V2sqC/qkz5APbhv38FrfXQKRhrvNmHB3IEPib0KdtzFwNgX
MF2u6tS47Wtl2aN1ip1UQVkrvRyPudmPgGhc55m10qCoRb7puppRjfoIpNHPoJr4
I+WHxiFUjMq5074c0EJT8nBP7tsA0GJILqvIF5gCxTGMt7FSV75dFpA3YjxhiCWL
owmPtiK7i66cGU1Z5pEczqYPWQxIZw3/g3+oUygkmP34ckdmdaN6HY3zSnUf8Wz6
jJSrWF5hptvWxs+fcQh6g/Zo4nr00UXHg2UnEtvunMZi7dUkKVqqHnONZY6qP43m
OCAPR3W4pmSFtSsGnAgeKmt4ee4Zz99ufijOa15VKFcDAOGYYu0vucciA9CV6QOs
0jycwuy7d8w6uF1QaLVxsipNBxi6aifR894yIk3wcAU/v+0oq2/9xOKNCz+laxUJ
FLR+FxMmXRmb2oxmMCt4+w5uCPqwlJs8gBvsLnEy2pY4z2mN0mZ8SrO5aFz7t3fY
RAIlM3Mn44150ACO5P/W1K4uQhDXEJ4stt8l8rCE5QbJqFFYu2opEwymLoeaM7YO
J+63yVXGA0BYg7A7pqc4KgSCq6jngp/l7fVL4tpdfUw8l94fgs3ld6xmI5kyqmcQ
536Nz2Ymj0rBlgAw28kQ4dfoJrit8nfQOh9OUOWNmejKxpk+BMCFNX7B6BKKUszW
A3aE7EiSuXa+wYNKOkTnNrR1A1idsVCggoxOgtLGG+xvLao/exMyjQrjZCm1NQ5x
3SKTyNB5sjInArAQXyZx+e10bBRg/8krcSC4amL7SzPAiGHIfScUDEDRBv/bcRFm
vzW2/QsY4SKBi5hPZBYR97Eu5iUIjd9Rt2K1/DPV9Yqkpv1MhOwfHHi7YbXYLi2D
U4iPtRQ3Hi8NhDVFeh9A5oS0iIMDzONO/j4ghA0Y2wOPzyBoIbPntWlD/mZmic+T
ZZy3bp6q3zRBCQA+vek44OJ+tAmqbLiFkOPUcB2jX4GtGSms2kN4xIkxeItaP/vG
wc2wyk4PbKZAWLxrjffLP2QJf9T8hPNXgQf9xI72Ek9QXWTGe19XEa/KZTiljC/Y
+tEmBP/F2FCRVXepXlfIjUMfe0Qu3iNircXqzGAsQ4DoMep7RqlOB+pcQQ/qfCZb
HBjk7WbsQ9HG7hkcwR6A+V58r+0z/4BJdkwB4zOIYuHhICR+5Q7MY8qj55VcNSbm
TRRKrknEqesfC93nbxqnY+4LJavF/MJOWa4EOOeCrDXubdBWfjiFCacG3ClE5fL4
ckmHRkYx5Cvh2Z0kLGTJjsCjloh4BngG+dPCT0tP1kubg76DG94xn+cqDMk6iIHv
+YbJNq6VpOloGQ4mt5buNLsR6a0pXhmbgcoEH4+MjQgEQCuOOItzDJ1IaWff4c8T
eAkUJXuofdk/Uvin23MWOPmpvQN+RmEmxWOVHAHGjR+SMUQx/A+1nV9hISAwAXMz
HTmggNq+ZmzGUl/Kq6jKLWj8LvlUwwM0tyUXsEEBJEf/9ZFkQvba30vTgemaYQLs
86wrHqGF+KsViUr4/5DbWZvkCkc84mdDeUmGXZ3PYlMHWcStIpizpMtRXRPREWCW
EeUQmsGN1mpQ6xLJ8n2mEWb4uTZjFFbWtRWSV7q/7MurubxECtAGEVFkJZEkF9xC
q2lG0cdjePG9V7qtwnxg20jXPKCIEwy9lHJFNhUuracJg0Q7hresNlocvvPUlFfw
yk3oqI79wfZ11hmB01PYmR6MZZEusli4h2hf4XS9UIbCsEdUbFNAPCtdsWtqaZMS
0R8nxwJ9QKeKt1XbG3Dx4DXNoTpNJFfGQpqzOXC3nfrsPXbTq+U2+NktiVjvUlEp
KvuHNH694D7wVZtwLSA+IezpU+iev7wrf3hXPaJD4iUGHDVjPtJP+hxwmBW7UPzn
LLO6hSA7AJ9LBS2JQcz8hw4FUI+wz+29ni1EXZN789eBXnXeHnK1yRSMnpjxuEgZ
/0iSpi8nV36oHz7NCUZ5ukByJaYdEgxeU9HFqDiN9uCHY4EjUy/xICtZbQ2LNTyg
8+AlrXuLN7ZtxLzL8RLplFQ4MOQ9N5HUBcjFYz/gAmeWbmDAWLhojiYlAEcvFe4e
2F5y+4BnMTig3S6HzO8k00QJ64VIhrgFA9ZMG62WJ4UbjPIDpxyE2RgfpOqPLyWi
ZaSZV3svUZVOiVNnMr5al1KnQHMywvMjSqpQ3XZ+3Fwrc0LHJCZbQSJTfq+V+1wb
EG3VFVz8wT2Ba3t2FzqoIaU+Smb0xrDgM9D+jdsBWeQ5McaEObW9hI4LscQo3GFZ
X7smFwN6ERA9g5Nl/oxYzp7WJ12Dj3ESxvi4AOzRKprwchecko59MWHHIDsBm0XM
1jLKnlzpmTmncEZsHFgINc94d89l5P9zRH2fHb7CkZR/M0cKZkOvyt+v2e4U5Pvx
4ocp1sh94XTXLkok7R/w+krlXiFmrZo2ViSdz4z1XAFioilDF2odKGsdVywCqBFN
MKY/2Xi2rwdHfzIX8MdYqeUjAZBGg+QDWm+BQKw55HFpwHFyDxf+Vken+JCjVJEr
vZyQscnyOzPpwt2jqWneH94mLnFBBXihggE3Zrd2cDh+AZgUlNRTJ5yBtT/BmIGc
3dbHTvQ86lj4CGtaUYCQOXc2SEFgBlnZzRk/oUUzZLVvpjOTY6noTHwo7RwK+OdS
e8ou52NlBJ9Gipe1DN9VeDJhiK++FWaZYmFcPZuvwmx6Z+BhAD+Vs0fMks+gFQ3P
7+eeiDq4EF7hx6OGAV1moyNZflSYGK6NPgS6l4Z7qkTyDfAJkc1ote1T4QBwJFNX
bJS19FIpOQoF0e44+ZSGRcdItUCPq4wmIPo6dukDAfMaoZP8gLca3VKsuZvTO0PA
H2MlEXdDDI5uNMllTFxOpk3kWK1hfIl/svBPlpBQvmiZNh5DCKkVOjXMVZydXsMc
HGX3x7iR8OhHJ59tjzkjJqJpKy9NGLlhwwfNMWQ2QYglmf1HShgAozfwyvGmHNMG
RJ41rvX3mkyxc2tBrgkJuu/oWCevwQu4qMtWsLmwhS8SwNWTkEIPgXL4SoKrRkQS
jTnuT5V4H8J23WOQOG/InphfbrSGHZ+mHKcCCXb5x5IjE536oWSiYKL2uUDY9NSD
F9Nn9+x6XloJB9Jn7zzT+jwasMShnO92vE5tJfsBvAKnKdQvEXekdRZ3n1rJWBwW
YPLAGo2AbkRvOqfWFIGU215xWYY2v48FjAKoKdAES/miLqtEH20tUthsN+MbRMvY
C/F9FMdegEdltOD6KlNV1nFmBnNOFR21Mh+76xzMYqlkAJA1VBg9iJZAMMWIrGiM
obmr0vm+HI1YACOFwU9jfl6zs1R6+TJ9+roTQEgqoK1dkcVozQlVOR6nkJyJ93oQ
CEcEpNmsKGAGA4RMJ+xlqyJ8BwpKGlqlamKn08kAdZ7lvJeJglB10JhPQAvDnR3c
gj4r1N5H0GkxRL/dYQzX3LgMxnQzsSFg/TGoSgTiFFvTm1R7qi+7wRmO+1IEWlTf
bMVzGEoGRurb1IYfy0JDP78zSMxHRqNvuqnsXzjMkrgQSJ3eH+zt9y1n8UEH0Bst
w7CF2fH/K3p/1p0/Zam/0XR7QpxPSJGaTWIB9XOGSB4xZmmJoR6Puq55+bkZ+6pB
M3aAt38MNn4S8M+LyDVdb7bu5gC2ks/4dMk/ca/rRLNHP7iZPmQ1hDPubQK7+7pR
vlTtc1AGyr9sRVk0RBDsBd9Q8BxtRjZp8KAoHROHgV6AH6OOEG1suN1v7NIFPqwO
akNQQ2LOoh0hinQLPdTMeSZ5ojNZFK/R6iCZMd+0ZEh26IeaKzEWHjL0xd7O9XOt
/flW7XIpHWM6mnwVE64sBgvKlsN4LRDk9T0zVAhiPQQfNn5Xta3v+TZFrnTinRbT
H4YKhDFy7/KQcKm6LtUQN1xADXfca91jjdKfbUQV8If27ZFPIBvBXmqJT5yMN8oO
cveC1bZb+s95pBM8ramNxU4pyr0zlBO9Q2soWP6Va2Lf7uFOao+DlfpLkrUfe0Cm
s9iDWxq4BdU4S+Ll4TkNawxZIgMnXaHiOxVVkPNYC8Gb6GmtMtEVNsMiiPIcUi/u
Lxh4GElZ7Pm9/PAAJ9Pox6wYZbwLGoWiDsG77oADzQVmWvwAT5hFIzw4nDjqkAbw
55GzWfBamfk7Zk8wpx3/vELN6/wNfiRynArIWQdFr2uYrDlfiq6J1lsQGI7xWNtt
Qq1tIRFN6/7MGR6QmS/OKSk5zJ9siJmd4/cBuf1wA88+vNGw1X1lS8n+tDYPsdWQ
Z1eL0o+hck3tKMCn0iNhCNkAdyN77YQjJjQAeY70Ni2KfXYJIN3PfwngQfvHMyDy
6zxhE5nwGQJZTr6eCSpJhAUy4+bzLL+NsMbtoz8+bDALU1x99kTRHMhMJjZ3cpJQ
y7aQBydwh3ZMUK9docpbuLrUmOP7yWry+h5hiWnwLKcqP8ON5iyCm4upnQoGSXJe
4omcnO4XHXlfdwW1+PS/ooqLN0z/vXH2rU+fSz+y3jMF03LWq+JyjswWVcyTvovQ
kJEoK/NLuMUbMK3IffICfHolgbfNGSI5XkC8vCYHWcUaz6WNlmb7yc7/c7YBO9zb
P2G9aHe23BpYxjJyX9ZANYh1fAtc9crjFSr2BSR8kBWzH0C2TRqRji3Ieyys0dl7
kO0atPcoRLeHRu58FnHh6QfPQl0tn6V8e+E+1Y2fUQ5FTaL5b7ypLus940NUMtZs
GluRzgrLB85wxC/yMBcVhmMyhD4lWIR61BwkVzGwA46QwDGu78qcTeYYPYNmJgMo
Q62mYDDCFb8fNhGTYo6WImxHpCW6mTQQhowk/UwJlUmaPkQtv3UZNoFN6uaWOVKw
apv4B24lM4ZtvYoszZsgF1NphPa5AlGjQ+D/m0VLztwzJbzkzGegwdn3Eeb5rpRC
FLry8a4m554CwUFKicttItRWlEChtMNKvLZ7ltTUJemIO7AmP69+28/hLqNsdrl1
eu71sLsWDUKZH+oE2FWfvQ5eummgEytjhEjhwEOBI/xa2CXjNJ/FR5csXj5EpPBd
Cu8R11C+m4SGarVTrj0dZtzF0OG2XQSG0qEwa1lORYXjhhNm9fUUmrHKBKfBzy86
rMcjlhQwHG5ynVxy/d4RCrJWYi+EWoRSyYqWfSeTdrHikFYdV/zltCBuB5QkTS0P
3rc4375PmNES8u5eGMcuwoaGJXArYsTyOJvymhobn7E9iQjaKpl67Zjl8iv98jUK
I1CR/UbAV3SXT0NUc3tJyakm0CHfmUQ8irL+sf7faqNPQJcKLtrpRQgh2EPBbc8n
DZwXvk151+Tuw2AoS7UvPSmpeN8cLhxBL+AAD9r/sum5QDANdoDoNxNA+bICben4
7v8UHL24yqNa1WUM/SVidTimcjwQWCMw5IxSFPgx2k34JQTxE0tIwHefiIYTo8dg
0pj07AvgVJTLNoQsAXPSyb6xj4t/z11tZZ6CiyxgDd/HPQyKr/vRafKF2ESGxmS6
DYn1/laVjj7nkYa8D5OS8bMcO3xGcUb9d+Mqb1+u39iLjs2KGeCaR82c1s+mZxkE
nhpdEFAhOGShOIu6ZD35SJTWmGJoUUCSuSuhprWSLKqVBFSCDM9qS8nEWJLY827Q
XqR9U9TGq6XrgO5J8+l3SD9RzwHIJBj61+Um2E4s/FOHQnYnVhRoMadCtKdNKsRU
vMz+B9u8rGA4FmpuocpIQrp9x+P7NL4tWstC9RrEWNQYMP5GQFTV6JHO1G+PjinF
aM2JrgFqH8K775/RGhztNuDsiFaK/FTqkXMYQo3hzmK+a9DnT0cBECm2uvakCz3P
mPwgRu+w57ma5YSVjVm+dBqiyUP4BzgGMQrR6Dq+HHKC4MQ+KK+5KHJHuuKsYpXw
QhFVKM0VyJqZ/FcwBbe0Iy/cEVMqp7ql7xnPvMm6XfysPH65vDadOjbPqWYX9Uqi
su5P599x1LWWGFx06iobe4Ojx4Tx0i8JiCjiMGu0B4xhjhXF3T6+L0lSVwQt/jck
irf0qMikZP/IAcEWJJuAE3qe0v1oWf1Ch5OXXpkwEmmdDkkhf1b+w2H8jXmgKFkO
ApNUrjpTO8zdqL69TdlBuAGZRyzKd6TQcVE3zbZEVp1YSm2wFRbf+Dhx81zPtok+
/I70aBdoNuNwSMoKwo4X9GfMNKXTKn9ystfwE6E1oJJI36D1hCFIsh7uPaRGKwcw
lEMtimTzmG6yw6k4Id7//9JWgBf3IsKbrZnXB5ETcYN/cuWxUZeFoUjRkXEh9ESf
JOq5YML9JHiL4v42E5RwzIYTB/vJic7UdAUafSpP649DcwODkW0BlPemoQBd4TUk
sztRbR54QoGWCLBZbpcHMq1E9VgEjgSbFt9VVUzN5Lh3QbDfofGNjx7HoBaqAotz
QLQvvgK6wwKEkMafdb8FeU7hbemn5HKDlMX0opLd04WBnB4+KTnNutS/2T2qCwZN
XTYggwQePALr3sS63fYJfrxTDhNxjAsy6IdQ1nHXkpUGvRrozjMVK75DujOfQRF/
RZCMN53j2KSQPX4j6IWGjQ7fKIDNpIi/B5Don7hy74vcf5trZS6rIEbKBgBX1DGv
sZk6rGDpq7gGCXAosWdxpK4tV20DSsintQNSuRm7QrmOhuIqElja4DLhNN9qLgKW
9zij6sughjt8ihvHlvFFTcee/mcFZhf3TQDQ6KRvolga3zyMf4gRb0rHN9YfbRry
zYJIDZVxj9Oo4fkPGT9tcnr35nwTa31HZkvpJE2iq2BN/+8pziSPg3ZUTLrj22AS
z5ZdjQm+oG6bo1IcwGr3Va9JAOTJqZtjUsTKczDW5Dt2SRe40cB0rBKo3fqD5ef0
SIhf7BxMrDvpm1P1o2Zyl2Zw+RDPJouf9yfpr+Kk3gWYnfqGKtINx+WWmMBe/VrL
FcHHbsgtSkck6wLtcMaS56p2pgFX/Rqc7hpsNdb7/OpuiMR44ZT1sU8t9JoQHWd/
LVtlXKtENw4VexE5JerIEqfzAblq38zXFIqz06ycFlkGwXFjQN1eKilyR6DbO+fL
8zfn0qaJscEfrBKMpCLyUZzJJyRiNTpBU9QGWlA7swZ8dMITzmQDfTwd3xx9z2Hx
0gskbUpHXEkZM9uBXYfUtLXE+P9BsAGobdDBsEtnirBi0Pyf3YjUwk19tM7FvLv8
sDh0ASDQlpACrCt/LghCKgMNgT1UEz6bQl7JhJDhHsSxAxQJmm/o/nQx/b2qYlZk
xVLQSv9B12TMjarzHWUpwhxNg3ngPHr/7YrvHB9378aD/ZdmPeg6HBVaZZFFaev+
yB4O9zUYO3ICqr9akTmxo0ZAASCYI4HJ6d2JEcr1jgvkSFjjrpUCEPmRY/g8tTzb
vWj0HccUhWhZFI8DKgc4jw4oXq8a9yllJxYcdKc3EfUeMOi7wkn9ovw5T912G119
fDbcGqvyu/EMK6BO+5GUK0hAMQl8QUZBRwtrMLwskGhCDcj1PZAS1cSIDSqOS/U6
bzWT1t7ITu88eiyBdLYaEI5/mE2EQnfqgvIsldU6dsQxluf/RerW85fdKImY/k6F
azO2RhzaUd8WUi6NKXQT6gnYND4oUhaDz86FY+Tw0YoixhaMM1o1//+WPveG3Ji1
kDPQlpA3Cq9nBILMSNrSNn+ZZ1XFfWUJdru3TXxfGOQj0OSwei8HsC95qxYOZ0Ny
e/fyfchD2oYliafgEFh/nvtGxOXts5ytl6uzVf1G9FdGC2PWxtGuGdQyXqqBVTwu
sB91USSK5hbZNfHDFH98oj54RE7UaieSeHOXsy4B9e3GX3K+fG0ZkPFaHyVUccog
+RT/xCzXAg4z5ugLbWTiQU6qKGyJiN4np6UmWJTfTH+GwIXvdFtVdPsOiRI4bc5A
CIgF9ga97JLtYnC/sJfqBLHoUV4dDysuDbLeEM/W6qeUKCNIIYRanztrhOFJ4K60
4P0A0TNzMvLoBYphbLw9gOiZF6bTKxGe3lCK4i81Vlh7ltPg9V8wGmQDJK0g+p4E
0znEaXn8r6UlKCwha+asdlRh9nht1/Yb94RPkk+MImt9Dxsol2X95zvVPAopSO+8
b4YKlhWthgVKICvjZ3KNbnVwDv740r0DA/mKkrFDWVY82lVzn4hjECxMaDzDEBVx
3ME7ZjYhAN0OO14lkd1y6YzzNIIhnrYjLMyR95UM2Bbz1+hOKZMb9hAmFkmcqo+e
1IrUnsDNiDAlPDvSr3Kqe8w0iOTOQZ/45pV3r643VLD8wdcjBJnzxTQcPpdDTC9H
+iYWIByKouZ0INmDsiGmxqHezzJqbGwaNbgr22o63qdo/azv8dX2HA7Gq0LZ26Lc
7DvCP6MhPErWcZITevcAUR+qQFQ4yiJ2h7bihkYz3tEnO1u5PXUvcOYIK+3AZpyO
8ZDaHGaOL1h/jPYvcZRcqZm6U8O4xUZ/0YGNsk+fB8tig6dKCLF+7MhUIzMG70kl
dsO2y25l+9GySMRVRPvMk6lA1a3dWeRFsmN4GoEqAEwy/e6PdofcKoPUKKOKE95I
VZaSYzVIcYcdTcd7PMubAiHYPVfbLP3zc2k1nud7rMqhxE8thZsNifnT6CgLXa8V
PNcTjXuG9pWvoNHGWwiHJRn2rQyIgwBRXOC/hv3UkKBKFE3FXLO2Ay7L/kqpJsJW
bHsVCJMMTUmV/GffmQZA3fbIQ85YskRfNO15+ySjljlQXcSN8DGTXDpHCV4dVqUH
m5x4k3ZYSo72i0X8KmMpntPlBaDbB+kqLAghCmJxwJ/gJWjTA66b6nPY5aadHqpl
MAihEnfRdRy/UD5nXcqE4/G4Zk4EjkNVQtaS/BlidazyEWxdtCowkb8k8SgNUoQy
6bOQmOcl3mxkadoeC28DZtP6nDPL+jIXiiBpUmFf6HwAO8La4IA03zVVZB5P35pq
NMdq4hKsObdoOuATfJEXU3rZ5SuLM4DfkblbnqlIfAxKzWIc6ilq0ps29Mvx0CxU
lJYc+w0hqp0McUR4BtdLM1tICUB98Il7SlDboguYApjLyE2iNz6es9CDPU0bKOXI
wMd/lMgG7K+psa3ZBQ+ojliDO6LrJs8AkMcc6kv/caGz5vel+kOgGirDcn64bfwz
Ef5GZ2+YJ8XdZkqgHbQ/KdtONLn8Qa6aqBj7n91NN7fOf8T/qwzMEkt1d5Y+YiBh
B48AP6Zx4sZahU5EOC7etQ==
`pragma protect end_protected
