// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KYeCLAfaMJFXNV2RHePg9k3psPQv0tFgV3lCdOP0Y+PoTe68H4CPFSgG+XzRGAkr
Q8g3sEp99tQ1mSgYcrW1oq7YWQahkaZuiLyYBzFiZxaYHraMTduryhA7UCaqXiTR
iacwkKQkOMp4Vh7OOMblqKQZKuRn4L9vbfwyq6s4h6o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15952)
1v/lWPkrSB1WK1H8yVYNTuVsLM6FSG6QAJYh1KvsUz3YduxRoYJ7hA5sRoCid2hW
8TzVTlYmoz37hMlFml6tg4TNUtMSfGA56fHtwiGtoLNPDenu0uZ2t/mbdcLWuuH9
RM1k/577+K06+dC+LZTnvpwLKTAH6x1k+5OkFR3uF1bgs9YumvEGi/IbcYY1uEL2
3dDP8IMPMxRCl0u3IC76mesAkIbGv/w7JGIfpfspYNzgeWcjVV8M/7iM10lNWXq4
KDbjKj0EYxbKXpAOBVIKVHTFHjG5Xxfv3FHMailvXH/nu2SaU38CvdYkKGBVG9eW
l5fX/Pm1eCkcpRNDgIiuN0ccIm+Qeb9Hmr/uIU/BZIybQ4tkrhT9wE8E263UTipQ
j4+IouPMvD9Gvc9kmx4ziyGNapX+clUYt8uwN939EzIlNfX0MlbGrWsXfYbDv8NZ
NqgTRpzgFC0SqcGQoSKkBMrpJs/4JFD/ARNGPyTt0qc1j5DSEE8cgzFHNAYQewaK
YlUjr1Pg8FQUUoefodsoAEHkRr7/6X0yzI0Ib67U+JU/f1FXcwnETiJ7tZdRXMts
KhspCXzHrbz5n0is3uX7/6tx1Y0M5vRVg+JDd8mvtzqKfpXaNts2q3jXG4/360nw
t03ZLgfoHSikRXE0qOwKgkoImTAo7i48qpF2c0ym6poBDNQTMsqzQeo8kVyvx/hE
awKMKBSNK0MLvGI9aZhLmMZOj/Kq3/9fDRZNYFKT6l0yNWce+ZrQ6oehGlNSVsmt
B/k/G33mG1AsF9vEvbo0M/fB2ZNtVmNlOsFTK0joIn1adbxMJy7CzfVrGo2mKKSv
ArF6zQrWb8q4BQK202AOseVuiVa/lNrZviFbqhP3XSV6vi69wnKaFUAFhtokmBTF
J9740cemzDwWWRpc1gh6sQ98W7Z4IXW3Dy4GOVkbQ9Q9qRCmjpHQBElSk4Bpy1IP
YK0KDvO9fDuFkZMaPB/x4YzpS6U5te/6Z7soMasdAFGS5myqRyJmqrjk/G+oNXwB
tTZWRMtAiTVe64L19m9CAd5ajxXihFY3Qo0vO4u7DJ7eJkw4r7zqj3eASFTbTUb7
ZhWz8FrDhmTCoXnGuH7qLKcg1dmcGySrhxKLzNyrbmhEMpzFKxhm8+7MfR7Azlqb
n+vt13F3KAfDxmQZmx4GGeLwFQ8pwOkvF/Jsf4gCfyQY2tvwQJNgjihZ6A70iUV+
DEU8Kv+4H555sWJSazzUT8x8W0aN7PMwnmYYrdPcOgDd6bSTPwx4ZJzh+aUBTAxB
2zNKxb4FlQuK6wo9ojp6zXBkf12igdJBNGkSlOvBtaNo0fi4eQTCm3wUR2qgRkNl
6/cVgZho16V4KfcauzwqFiUtqf5AW7BVG/yyRvUfiR5skJkJgUFvORPLeHrp/16U
2uuE6QWJ3/IxqBXwPtsDACwMo1W06VCxy1qPH5tzcqxheNCfLDmouWYE10Zl7lSk
4ZlsBM3EuR5Bar6g3PLk43ojHH5J2KxzXcDGqggMtVBjnxOlYa5F5YkIFeWWorQV
7tDNx/UXLm6WOiaDACIhxplllBFqvNsxAJiQNR1hZXR/bhiOonAJMIP2baxW6Na4
gDmisLGURj+C+DzsbTGMwW+aQI9YN4iNdpigz+IUH5SLTA1b5Ye3hGtsOndyHf7n
SoB54ekaTPxdKdLXwJ/yFM+3GKcuy7uNvJNbq6uAd/wMzR4s3LAXRe4AhFjvRVnl
vDserzUb3MHOSSjw0ZbpL2HQ4M08ufgfk+VIu4RAklOjwwcZ7ftcncy3T2TWc5+5
N4L710oDUKG0/QEV6IiAbtrqOS3j2Gd7pXSVb7C5ZnD4v0Eus8QV3YMwQm/2fzBq
DsbL2bswAXdqGEiOqBebnuHo5capWuqQHMnxpViEWE5M++KV7NtF9nxpCz2gMu04
gBYcRrgdxTSRVaBxNY4VMt2HTpxyTj4wAqrcFizFKwjkPNWioLUR/cb2CnG/w6Rf
xyQCoGPhRbEDlh2NbhwotK4K+W+4hxFCDgckhmdDylJZHAOfRt5OMurolIPUloHu
6o1XMJDP2vHur0jTFokKcy4HbxOmP9Y8Z9KOaI8CRs8wpjUrbPfeBuCB17qjl30E
Jzslquyr5eS8NBqdjuNmdWsWuRAE+8w0JeOXhG4qP9QuzeArK3AfrvWti4s5Qsth
hQP59IjCrPAmXgA2tPDiyAiE4RN8daE1b1c/Frxl5D9YL4X6JLxlUnKoIiMceQCU
eSkmJy8W9OFpjJt14DF9ZLNyODxKL+c+Cgh1cSMG2aCDufsf8clv8vbOvF3Lm4B+
7Eexum8mHeROxR2WHUppQqwjqdlLyZbRA1oDtRGexgjV2R9f+O+ErqV9NRHPNsDA
WRhhPvN29WhT0lk+BD3jC0JoVIvmF7YJ4w3ex5WtpZa6QFxA8JLh4Z0b9fXJjTB9
16756WCvfhRRB28IP1mhJAOYjgZFBDavMRyfmQMoO6iWaU/1eaocpSAzT3ny8Kqb
g//QoyWv1vVcT/kei+O1y2dQUsfRafVoaEH6G+llXLo6/xLWzRzq+ffPXOtNHKLY
wvuTXy+b1ocIvOdCfBrZgOpdc70cl8hNgMJzjY16kkJnvsXhwrLn/JcYvi17X77U
COFMOffYnCPh/Gq9vxaCc8aO2DnZMLYdI2KWpTQhlD8TxUuW5ulRQYsLy0aDwmlJ
9HkxML2r76ylvQXovTw2TN4IwFGnwgXVZ/NJpJ4z1mPy3bf96SDFfFtC5buwZCV3
SI61RZXg64W9gxHzX8TkURDDlR/Mo6O35TNsAQFxJ92kgEJE91/BBgMKFPU0eX2F
oTLvp5Ew6eyw6HJo6BV9mmOAlQldpSdTZHs33+vpEtgrQbfAFLGxJm8uIQeoSxE6
Ml5e4w8iscHKUXi3MQD8mbeHWvAqt7L8Onn3oHluOD5oOrXPcYWUHO+5ETrh7hGN
tkDOQIf4OvXBQXYnghiQMD1eRNBIOz19BMMbmGIGmXc0LLfvK/iHd16AnNRmAblt
y8CyUmtJXdzjthb3QCWsP6I099RKJbCxlF6DVclHnV3j6v8+ozpWUpIUGqU+XaYb
l89thgWXhiWxbzesvWVQa+2cfuJTX93IqEZzW28dmsd/0Fq40ypxXfaEsi49jQDd
/nT/mtubp2KqXa2wqaW6j9OYM44r/uhP0KBkXo/7aG36I5oQ1AtiQDr2zFrjg11p
Q/xu1HXx91956Af8yQvDN0SMmo2vW8x7xCYNaowYrKIMBaKOKaTObggMdh5ORkGD
UL2y91uall8OFbwnxomsD2dW8AhbfknTCEATieRBqZv8N4lVwKh47tyWP48VgYe/
Qkp3Y281tFttban41npTBqlqYTgsYDfP7ylM1Br8M7arzKY+apiJx+YxwVU2NAnf
BzDPXe5VSBbM2N0dH+cGvU3WIhwJAzg7nGROjWoH1lIc7K8b/3MO8U3hRrknBgkB
ExAitKI8U/s9wq22SyNFa6JcLsblgWKPCKXDhIo1qCOf66LRcIPgAiBh4AGQfN15
Yo8M6/M5xegj94cTpq4BC0TFKpjPvbnPYJRld6zyA/scUfZAmLmVF5Q6ZFcMKvcn
rN5ClErCSw5gF4KT/e8uD7Q07cgOywSQBl63B9lfw5CtyGXsTkxKYdp7bTtKfFIU
u1bNlwXz8EPe8h8cy1NJt9AxiSSUat6VB9JYhp0BJrkP8LWCwSwb0W7uqP0KNK13
xRV1Jq7TjYruLs54/0eLxfTdEZSF5xJ2/4XHhkZd2+vfuCpxV0PYvS5hfNpI/Aad
TgjlZSKf2m1X1sfkgCyxUIOaPnL4BgtlEmcQwBuJcloNzHeiHB+0lsHIr6hGdx1Y
S56XgZbnk8G4QFj650j/+VKvT0L4eGZnCFEslmSs/pI7T684cq1QrISS4mQlK4UV
TM1rKEVP1HqYhOEtCdK3mmxcQrbJmKaqiJtsR3IvFJMmZkLlJWiFxbNdwK6s1YaS
+FGvSGHeYbUawrbY+jn2xpL6UW2V6Z+5RRuhpHNnkOnrk/q+0ZoO6QyzYDtX6KyC
BCJrvjQkuHKcBQxofSzv0gYQ8LIrk8G9gPBeiYQph4QKPXsKtGJnyW+bIYfr54jZ
vBHxo1hIEfz0p7oGn8o4gLD+AThcQH3oEuW68m3jIWTC6tTwYFpzCxDJgth0yuIK
GDhyrZq77Bs5WGwNwlWJyICsWGe6SWswhtF04yXrE53pkAocpl1H5qfc517gD+QG
h9gibE/3t5tVMhMmegqmBm2QUjyX0LSwvkEVMPLlzjGB1QRbgdPYJxAYvAVouZ2r
zvUKkFKzMwmVo/TDJvbwOz5XaFZdoZN2fQ+W//qHmgbMO1Hb+8CcV/rZO/FX7T1N
aqxF6YcAcPDftuZ9ADRx+IBw9zLI8kmHCwObpnVX0WcHoapAYYDvZkGl27MOW3Y1
AJRY1P7VUO6bAtPLhGLo3FgDnsKJjL75pcxJbvhdbShvqRlN7covkCDzqfGSl3XL
yazRSjc9PJLB2+QrzpyueS83H540taAEjiAkC3sMMSiVyf7tVmq1LRmrdu30BcTY
S3VzI56ly9pe5hqwp8VUMklCIaRhxdvO9xYWb3eoDI+3UpYhPWFKQfk6Q1/91lVK
azgdylwoD/4BbLL+WJZD5uPW/CcDqavrkxLaG8KQQMBMUGAWcgqieqb1WYkA8v7R
Vblc0S9PZEc0mYysJWjvojbtBx7ZU5Z+aaZ45mNo1k6N5lCUABAAqd6lgEnxDNqu
wLA7ZK06aFaJV7cisdP6m8qjh/aL1dq2pRHHYFgX+SZd8VYWIX5q9gdDHgiv4gXS
6ZHty39J2QRPilfcrU3vNfBHpXRl0uj2N2n7b787khDFPSIbgsMcFCVPGs3Zb1Ql
yopw84i3XoINI6lXDG1DmOpSqqeN3OtlmDMhyBBHu9j0l9MQjlHmFNarkKHZiuoI
xfgix6gzhNyvVQzg84dmHZ07uEMbXN+T+ZuSSIb4DJA8biqQAxlPmnFPiZ1SMNra
XCXxUQ+i6I5It3ZsLoUdV1AAyWUEyyIoP3sNidx6Bpc34EiKjJJkHUoBUPNoH0Al
ExvcgcvVauR7yYfzS5WrX5eyx1j4BHxR3uHk4vseLT2yQp+RgW9QH+NFhDIrH+tV
zY9LNSn2dBWo+U+Etz2lu7AwY019dQRn5gsRg7BNmvxq4VfQCxOxxg7z5tzCEynm
hzQGLeXE79kyKfCcWgenlvhLK9kqBool2BkUVWZ3QQ9BhbHmgBaPFEg90H62t34R
AP/UALyyRZ4+eVwnqlYmsGL2T2bjPFCOBEvb5zLEsM6fiJBbZBM6PQIkTFhML/zO
CkniSkwf6ao4HkT6MI/H39cqx+4kbKoo6v8CzvE6QPc66oAwg9Y4qJN8d1KKi5dA
75KFHLmpN+wxKeFAAf0WLUtRDB9mfvPpORP2T/KhXmu6cVvpUorFgJPGIw7sA3q+
1/Ng3NWdQvIWCgBEjOHzy9BtbVjkar0FvwMP5j+tfWQUTCrnQLME8V/5oyTpIW+N
ESJZgFwbqUdn6Fh6JqswUJKfPsadALeNy86RcYCC8hDiG66adg+hezNOV8jUmw3H
UzdI5/OrzcbC6GdPhw/567yfPMpHAlYoeaUKpzTBuXWCncDldhtFWx5Or5MOo+Ai
m1RWn99kHz88IKFqH7yIqzihpCO+UaEDnQfL7O7zVFj1DRuuBXR0gnOwWcPqnCIX
DgkV1ZxLwTJ+IvhOBkNoext7VyDfquB7WzF3RFuFb5ox0DETEOj5tscG35GlrklB
K4NwFMtneGqNqMU542xwLLSvC4BqScON1lqofwIFQkYxWjuMcQK6tNS5tbP1vq5R
5mfkGpV5rmzLISQ95qFyQJYZ5UDGeZND8DvAXQRmne2bxiKu6hhx6EN5tBkTs+7d
9mYpYeKRWGO+kgvfPpfA7pamnDm/u2V/jHs7NiafPGd41uuCmdooJ/wqvyz1ed8w
nGNkpNEdZ7beD29xtTP1q17xok8CXyMnU2wNLO3NChK82fFKtJLPN+ZjYfftykWZ
LoD7ud5jzS9btjVMaPQDcz2siT0Rl38/MJAhiOexT3Ty4Zzi2dNNPT9hHnvTYe4J
dYM81IpMY1UoFkrP0xM5W9ZtEpuNt7sbi5Asr8KNjHcUlAf5awGcoFLj+WBQ48M8
lWMoAdTRxDswelsGxKh6NgXgFHa5deTFGbG+YCpGqZjr5Zc4aBfTIZzDKQSBH6pe
xO3dPidVd5mnGAcBgJ2/3P0VLqpHuB3vlTosIZf5CV4G0pu7YGa8J/+Ot7zH/w6M
a/aC6rcMFXs277QdX51GuL6sHAwHlIz7rYLXRZ666Kiwr/OLNRGYnEPzEk8FYzQ7
AGctXdkR4utM9lnFNSjHyhGZVHnl+JtMoBCpb7NDRiemHA+nagV7wDMYg4d8SbMP
LJIjNXBJlnl0tCYrzW2Iej38cPelur4fBW1nT6rnGf3/9/GD491Mavr8KE3j5haG
mYI9UvuPhYgX/u4+pZsfKd0HrclJ6kNru0rwo1xU9y/N9DlKMU48OIy28NMljx7T
c0n3nBsyAxhePjH79lunjHrRtNdlgnrqv9lfb/jUoSXZPcGSzGzsmXLoBgz1DNny
VjOzPCfaldtxLObryKUSCTJDZ1d17VEWXtN6vzWU8c1s2v3cCGJplsQfkTeUcpIa
FvpBIrNL65iYFkgC5ZUjGyACG3fNm8qL/Qz4K/lFxLpM83Hqe3gF6lQ5YwnJ1S88
D9Gw5J1TkHLI0GGngh1y9hTlLQmPKVLjUR7l/ps/lWS+WUZuKwvGZoPTBmUofsyY
2YXa8BKz8NxPAMV6ljpWv8HogdX3/hTJ0R7/rKavWaakaTVS9a/4nOPkUViNfTTI
Hq3g9rxwyD3WAN2miPp41ni2UJ2eh9IDGEy5PImPhSXQSyaoEpXa8fjVKRZSfsyG
7ZVkSKQj+4uUT+Cs5fjtVQj1kewbMu1cz0TdrCaPFvsENc0tT4savQgC23aleU5D
yoDylrNt9Dl4G5p74q7MHtRbY1OWjiKTB7Vkz6FDm6dTV0GXs1X7J5wu8AD3X0CX
sjsvho0SElQ4Ji/gtS+4PqJnb8EfzOBdXnGDz7CiwUgm3DFspQ7rYS/LNzdnznCo
uOoZiJBDmhBXAk/w36OCe+5mNXueVmgrTjsNMhhUaGZ5StIO2NIOg52bddxXbhNX
qGH08TS8O/6R/4pFs7MAWtkH4I4FthLjXqqFU/WFw1P4RkIImkMyBu6sjTXyRdmd
x33SN3k6AnoR0C5wdM9+LQQPXIJK7PBEBI91/rqJ2bfkT420VP0uFx82k7MB4+MK
7zkHUnnGJN1Q80AWoK2w4mj1eIvV3ModPHFHgMOqtej68HhHSe4BW+pBpVXPW6Lt
SVR/IMTeC+DrBQzCY5NGmpj4cIBMTXrE8GBlVvDllaDuYUSROR9A/3QfoKaSwswI
g8uUJyBLiFlj95JhpobLrbUJbZyxC+DzqIQEtBJ6241XYCXzDHTu7rQV9HVJtN5Z
vlWuzZkCgv0ntjNCc0414MvMj5yUAG2YoAxhoNxoxHwdAtx7ULXZAIu89GR2+l9N
yAioTEoU2KOw6/cbrCWTsQYtg70SA6hDkRFNoa9nI8E0EkkR0hHdKMZB6BFsd9Rz
41JmBGC/ESEhoxb/fiXICMk5T5g7sC3G+lVPsK1l5Tuwtw77MXCO1C3wxdPqtMdH
6hXevGkpvdL6+o1aGzS4wVO6NueEboVoJMZRabUpsDHssZ9UjmLm1OkTwYn1WE4B
fVx223WKhEiKI8JXNPjzr26egvDNiL5WnXSqqL4Ohe0oKYwz9R5Dt094XnAn8co7
hsHIt434YBv8Ywdsi56CdMiunJJcn8XpWKL25xSDxClOLV9Kcm6aDTzmxWVlwH+v
C/6ybCHZQjAUdZkVZvoRYKwMA0k5llXXrG2ClGiW3VFnCZ7iHvkptmoWTwd9aXKB
uYkUgFozqFE/gbiCURgRCxaKPzCRhxA2W4StEEUuYXdTAazdlbfUIv6w7ZImmmRz
HFoSFC7C1aC4EZI5vRQEjcJy1zlznpye065SJYX+XCWxn4qGwOCq/aA0o8yGjJKp
KUjNUlpEJ2UmvEhnjIB99K6S0DsOE3ikHiwE4XcJgQdhIOyRIJV5npgvbj4OZ54l
QLblqqyYKHBtr7IVjEkR3ARghdGX11gifPx2SfwMjvAxufDr1kyVXCYREtBYbA6b
1CwBs/Ow0IhS/6dXUEEvEOrLVMTMYPfQh/aJbaAbwoBamFmh6naIrM5sS0iET7nK
1xIUEXJkcj6DZ1Q18kxtQEAiYpHntXVyJHgRKzVYJviVSi7kglNRh3SHsxf7NcSC
w+sTXHzPeJa38KKyOEBPrnc8Vu2haUOcKk/4nrCfW0FLmNoETjhgJRxPA9U59xOd
IdNniM7ZcK/JlfsJcU3MswNr5ZJBsX9ec7d86tlWwZdOhqS6OVp00ztVrM1cFEcX
yusWvWYhOQ4NJY0OrE9x4pVQsbgIiOVqOZtkYzKAmZDBObyHuanSVVPES13jVDy8
2Wqb/bekJAil0pM1oBsGMeKcl69Onzs0JlpgBaDBggX4PqAcAroATeOkoILtacKL
B0LH4bCVxZbjOJe6Sk8UFMZCeDqY5mn7EHoqRuc9okTEC0Ynv1B9DYnjcWgoERIi
tT/Ngjs/4nod2Kz8s1OE+2GlAv8EGKE1cVHztvidF+KK+LP+PximkL/L99vmy6Pr
398aCoR36O8zeyU+Pubj01KQZpTTyNa88huLY6p/avF59TJkWu79t07o5Fix2XpA
MSwbP0l9ub26Lyz/oZscSLJigdSBd8G38xDPzwx0bmAp7okDuppDqhDVf4W9gzTS
41PQF1vstwPPY1K1iJzmAr2SBR0iTk/p5GxockSzBex9mj1wvx13pNedrs558bBw
90NdzJJeWvc/YeWntLZR46TymdKVMOrxyyZ+f+Ok1Ziwwq7pQRa9oMyXDb7BmdE4
T3Uy+Clfwie32q97JA40/PsmlEBMGl38Y+s8NbuYP/0H3xgD4LnTTGfkXXPISLPr
vUAs6Zx/x2K33mXdlDPdl/LI7UlohZMANnNBJGj4/eSemBunS8/EQG3vvX/glzQ0
ZO8G5C8jIJzojogG+51L9UxJ5ie491HpL7I0EGMBy5WOBuWBpGF0vykpr7ncCnL9
m1eebMR0Epl6EP9G1oehjFDeOHIQGw99QwsI9r6FtbntThdzRCejml3c6aRcNbM2
j+3hpr3KV2/0/GABx5iR8HTU0wQjdLqgDV2gS/3kyYiu9TEaFWoKTGuxO0+YWe4J
h5YBlj9bYFsPtaFq1yuKmx2iNBD6nDmRIwyCm4QZ12a+FFNezj9W1doUFzDFN5pG
bzY8fG8gonGFntnUsLbQrHuJTv2j2GXHT/OhMSRANnU9q4ol9lXg9jx8HfexW+8I
vuk5mN0WyifC4N20m3v4wf3YrY7udEdmYNimNrQ7qLHAoaE7QMKvv8oAZGhLjinN
+lACjDHTdq9YnZM0xLrFDnlqy7fmlWFY82LKtU6JwTuCcPVBJIKZiKP920nGeEs4
1WPAr/39OqKs3BMa0UUTALVWUhkStxlibKqPrrJGTe66oPk1TC1dP/bmorGYXLgP
YlZWyNai13J7LApMrB0GxuP+5Bwh6nVhpQxeiCauwPEfN7TdLQKZyVIcx5SiAkDe
5KF/G+zNn79tYB380M9qP/xgQLjYr3tAD1UsD63GMhbLo1nM0a87gG9Ix+7+Kqdl
E3EDv6I/tcU03Q2EuBv04zCopwtlD1xQzri5ZKExWOETw6RUp7GO2b3SWbZQ8oIK
W1S2hYDjjn3QAs1gpo6bZgccMXgKRVoCWwuTG9hWjaHuUSipsWsOgTvBX9YTe90W
fb1/62vbZ8Dm41OPcDwShDzyhpCpKWesrtXSBfFf0ENdfCEVqbp8o1JBUY5xTJFp
pw5tV/kOJUt75HqXssI3tz2Xbto1NpiYHJ26/f9xWuPDEylpfG+3f53xgamqJk5k
fLgx2zWUNtG4qtM0GZiu+siPiUzPPFTfrKlrbA7Z32iOaW0cxFtvkIRfBpmaWmQS
4CLRNJHQ+C5Z7tRqLpGzOraOdOnK7BfZHnh+Ly7zjgHRcZ7Ms3Hew38GmPcmr2BL
sHCeh0KDXVcXYeexxdXWSLhqay+8FgYRFLpYErJSio/fkM17y/lBEHBLwyYIbq7k
Gt3Xfj0Haj49T8NbCuGzTXvKdlMbS0ukwRrojt436ng97BnOTzjiBHWK3Bxrm72N
GjASrGKUBYLR5g8ydx2W2xOqfjC9+41HiqNd976A1fn3wQUqGCLjcW2zqeAde1jB
UdAVM5Eg2/EyY08ZFz0/okBRmPrv0H8SGVdftGq493KRrTRcdyXXVCvvMgbaLp8N
3nLhkx5hVC9WsVZ0SkwesIrpF+3VUmB7LoI7t16NNNj6wpGb4jOHsUJjYiR6mL5S
eXeUrJENtKsceSnDbqxG3419r0XgW3c3WjwotNxklENP/GOLtKn/L5Gx2epRHwKv
PsnJI3UMkBtNfxtCwwoTBcl++A4PsL/LoO9ZjiJzIcoFf9mJMNgv6zecgmTBHJvq
eRTyWL4jY+JvaxdcS7w7yB2lmZVcBzGWQl+sgkHtMYd22CqUuRIhin3BL7eheT7K
mFnerpsX2OVLVLjrvPKJGm1PC+u74xGawlQb3X+DC6/AqXRXorral3TiRponjvFY
aOvySCSDo5iJ64+4JIzdoJ2j1UVP+YohU1YpUBJkXbAvhbMg3WTbURQzGRwXDQm+
WZmym1JY0SCpaSD9h5902wDmpoKPt2ih/mrYDJhsHBoHgVZAsA6pa1eoB4TVEfoI
zuenu8dkS3LDRC2t+XnQpFJrRxvIIJ8I3gwXgisScPtJaQuOZ69zqavkOA3blPqD
bEZYv2Gpunj2v5KHQSHAZamUhWxm2m8DZi3Qb9TSPuo1yUB/u3JO5pPQrEaNbxUI
n4gmbneJhtDEtWRIomyUl6EnIQnmHfOg4qdZtAxU+IBEKPJZBijrs5hp9pt6OBuE
0rnspcajj9YdI/LmKbc+BsbPP8hHTo84bb7Alcb5CW5KEJQ7Ib9gWNKvcQjmmMVH
dIdjIxpPQY8qG7QqJ8qwvC+VEJK44+JTeklW+nA7L+kAHpcKT9olfVbZbfoUbAjA
hrkeAAJo1yQp9EF5bJpHX1I6Expbh4Vo5Iu+K9Gv7sHVqlAuZQ71b4ZGsYgZ81ot
ClPgoDBlgphpboNOUYNo02wo38SLIDyBs3Yi3wdkQqAh4nPMibuBvpc5c+LHcuop
mQ5GXN5zozNraruyqdzhj7o/fZO/egUWbeqghCrYhf7njAqaNRqBImU9b0ZicvGg
FJ7DKOZC7di1AYnnkIg1gFmGgDxgtRXl976Q1V8F0JKsxiUqa3Oiq7vxq6/mmZGN
bhfOBBq7thH4OTbevqpFuowts9t6keb3S/DWZQBBqvhWGmuhPv+7O+TxheX0Gdyb
vJ/vBGivYwt8pxl2UIs9fLNR48ahG/+bguD/7yRjH7ci/Kgzmypze4dhh7haoxQ4
YifwEVnxIP76EWyQKP/57WanZC+fO15j7VzpgiTM0hO3rxbimjwnBeUeSStzPxjz
XHkS9ptE/Jcl9QF8yj1TtXOj8XbhbwvqYvVgtc2QWlMbAnjjC086rNo9WVJu97l1
fGP38YUgB3HqQDLmgkl2DnC1GxeJxqOzxehR0eWWZAXWUB6baCvBt1OWHnGq4kg7
czRyK9M1m22kA6vwgRcrGvsZWBh+Y/MRvyaqNZlLBEPDZpeVZlMmAmRnQsoyU6AG
ZO+YD/KIdTh735lO7wIivEpGm783gY4b3E3n5FisgIP4Qr6lhx4CkpaFi82j4RwS
cb+FtBrJh8BhkXOkIxUxgrChyBPfWVWsOO0r5/Vss2kI4Sl/fPLMYWd+KRIxcqG7
88C2UEHX6FDCyS5pVXTeQTYTmTa38fNr0lbNhtD2nqAfWh6yxaLXGHS/Ffuf80WZ
A/vnJJuydN9feOZBxRavhAX1OCb7OGP2l4P6Ntur7/A45qEHhTqsNwmg0NGgp9pu
0kQ/O5R5uCKWjYPfon6RwYo9WwUZwXN5DYNR/JW7y80a9YcAp8j1kME1sieP0TUI
LvmWFc+wB6RAuN/dCJ8aUADO8HCnrwNFNg16X6E19fmEeL9PfV5aD2R5q2UjrGhi
ZVy8fPJInCwhPTwmNNu3Rl501/MhzSn72kKfbIaIi7KTUPJuF8wPP3LP5RZmZ6lg
Tz/eEiRUiM6pbCZvDJAx+9F7sWSJiKWWLS5/0fGLLORIzr58d0FxgB/YWMCpEbOl
5/chDw/XTaVIfzrUfGPaK2D42wXQPa8Lt6u30ujdF52buIrfIrWsnQc7joIjBMgy
e7wtpC/1HC/sl04AEuoc1z2Yh07LkgHvvtZPhyvLhejGiypM0/d30CUeSleIANoa
cPQaH5kEEacos67UIp6mnqahmcS2rfYdVIuwRNmGK2Fbx3d7kXj9J5MlczmKPRcP
b8BGZJc+GJVWokBwlPgvW6HfP+dTlRUMTj8gU7id59nPifUYrtGAEXDd2bgqSVr0
JY7ozzzUStCJ3f8EIc+bZdsNpzgtLKigMl/fjm3lW1rNW6ofi3//MdZ6miCa8mhl
jcRkUWnb4oKyy9O8dLfy/Cs415IYgqVIdzdINOiEEvw2ATwDjFHEiaXTJJgo3NUE
EFSmMcNwx4/TEIv5ZcFuog49F3pmO2v2m8cyxyODTAMYIG9WTrZX1lAog2SiXv8G
T6qkWGjlUclMJyzaSS5eIgTluETv7v4fWL3+RgTJuDZILW1psfxNqK2NKXF9bEYF
XnG0oGjEIsjq501eKDFmJTTR8Ax5X3F6Dw4taxwBG3vJwREPgGfK+i3WxxPEyMpq
s7xpomuRB0G99h6MZ2956p666dSbZ2camWZeyNcDqtzmptp1UYgR94cq8abEdrs3
h0eupopnPFvrewYoaQ6IrAPI6HZv1rT/Sh8oqFAxiNMgwh4Q/3ukFcLi9RMUkba7
EFBMVOmM0hmTGPFQJoSR4Il8OVB05q7rAu+vGzBeyP1qDgPvWl1tVLdtHUnTptzI
3aQy4pwSvNSY8uJPfxRtNJe1QWJBe4qWk4P0NMOF/kAFMQ5VqyLYw8fYhkU5Uzf+
xRDgYK3m96lwizThoH2DHw5H+0VobZcYmUk20aNe5kFvJ3+4+LCo3L2vEmcujrN2
osIYW8xfvtd6orzWBvlOFHQEWmqZOuVz/4KR3neyX+C4295ygTjLd+z20cqTQ+Xq
R2xBpR5VON3kskQnCW7BXCubh+tlP7J0OYu86svmNYe+Q8Wqs9XsQZ1yeN+K1jh7
eWVeMRQsczSY6RF9iVlpV8Me5yxgElylGjEcP5Sdu2LAz+17DIFD2s377pKyrCN5
KEbIl0C8hsfLZYyXUS//qL5FoeTiMY4/oW4v0LJwYeD3Tm8R38nWVVWuGWG7F+8i
0HSffmP5j2S8ZYs6b2SJ6KrKmnsxrsACT/oLB9b60Lq8pHv64b425DAPjfeqljzx
LJIPV12HGZ8O9GTdjzxllV/sXrb3+Aoo0Pkjtd4KSPEQ0qXsJDtT0143oUR9jkg6
E/BJ6+4EVoCgsg9V2Wc7FOcOF6Mjq5L84CvaEYgSL5w+XFLD8e+h01F8My7YMzYX
FzwZLbN1UzI34hDIeey7OBuldRuL7Pb7AXGxCoNE0QZAG4dIsS46W7+HJNptj8oW
H0KasoQzYjlad944ET0nRqyW59iSCOzEnjRozScurfCUEoOMzbgQHPO1NLvsauhV
0Y1SU+g3TXsWjRI1uiV4GqzLx9RGFiIVakVu2s6nUgVtRadiqwuh3MpvV6sURdxI
ZK7E6v7440s4tXE6IuDJF6Oa0WuNizYoK0ouWLJHRaQ+1RDdoy3YLtmGLapZdw7+
7tL7xFLMlV3X6Kitz3gN/43ZeIoc1fxg3uyJKXmdgaKByJsVNWhIsIeEbMUo2Zts
86KHlVafwOAvH+PUywe4L2BmffZn9OzNWhUopny3VM3Q+VSyc+ReMBKfa547wjru
j71fklp1JCNVaXdWyfxV70qY7ewKV/d4lAO3hex9WWgXvCn0c1ACzzNoIEdH+MpR
bBKu1qNnBqX99HaApY3cSGRfYGQwBM6nWIecqhF4Hbfpa1WQ7o8BEtqiOP3DLt3h
UyBK0bAdu770TeWwOQNo5KTG6xAnoSG2dlI4jmVw7GfVVfyjDLvND6b44ngKfs94
Z8yF1bZRyBDsF/AAQVWaOsifLpdMYDxxnpdzB8ZNHFvc0xtz874YLTz90Tza/+42
Y77GVPsPlpYYNngvNGjVUC5jyJA2t/8Dr8/PRCnRO8TdRikcqR5G64p1ln2WrKMS
k+KWGFa0lfM1QQoiKrcY0CqTf2Wh3KcN7jhMl8BbtenGULsDhuZijFneMPPD5wFE
Ozd0DoHWQSeJlSRbMkOUujsDqq08EUTQT5NSjt6WuTeRRlpYvc3//xo9zCJn4aCg
r2RlvanIm7ghKQdd2ljuuLnS+PfiOjgSGU2jUaHyxIc9w7VYcdUVEOPTH4Vh0zE/
Pxr3U+YjEmay1Dp6SnTsFvgxPFLjJMZuJizzYTMZYXu0R3cLzsuViwY02Hx+87ft
36/nMBlummt4aPjROIfKQ0HE3McsT+kNW7JVKx9C8xMxPbcJLz2xwocaqq9hw7iR
B30oicEdNFcLWDoaUvNHgIcVWEzoHPZE6vDlku4LP3d6A4Z0L/9IUPL4XcNlP9J0
ONwGBm6ueBz0Xgk292FazKHfC3cbLza+ka0L0nShES/JTFPKAHtPaNXbZCWyc+fm
KBetz3Qy0CIGyyaE27CpVTq1PL9KaBKaum3VyymNM7yMV2mPjjpNCNvGsKN9P3tT
XRVGKs22R9UDA+OMYDZtODx1qVVnpS8HTSSC1fYiQAOhqovbBbXbtoWn+Os1d7fH
oj/+La7KuEXVw63IOj/NdLVEPbsuMT+vv09AyHE/gwLONhCGOXBK9pCh01Pu/iuy
OPj6D8kLIeAWHDqrtrL5mz20bjnvqkcadF3J35hVtfh+u1QqVRN3kmhsRdKV8DSM
WzlC8DRGeSQru4e1MGYb3Sbh3ak4AZvGtadJpb4MNRG4SAymZWZ6wiuxpo6p/GQH
vrvVCfdcqSV1x2sJ6LBP9OqLRYz14YuniHf7kkCsrfgfObAryLyXqdnPWXJY35gt
4iQ8Ss05Pxoq2nUBV9EoWCeORsoHcIaZrZrGRi8S31NQLZKDDFJpJFQ1nvla9f2r
JdNhk64iqyWYS39FGcWk2YGWVwGlgQOvncDB/kc9Y+IOVNjSD5KRaPQDScTwYhvl
W0xiSF0Nt6UKFCWHpxZPpqOwVCrAw5mz5AfmQXpA0s81Cm5Xp5Ky3Rpuyt5aabjf
z8XIgH3FQ11xmlXkILG+xDr7SN0I4Kyzdc+UWpu/p8Tp8aG/XW3tZ/uYWC7xIVXT
ZZhtdag5rzEbhRv8bbudKJjYmssCo1kQWzsfiEN6uv0C3f54l1TsMg4pj4qOVhl+
j/QaPIYFOKWWkG+/KEeOn+n+du1FQF5EAhaZ39BAVWkdLAWizBALBdGS6SpYIvpT
5Il1jAjMhzMREroJmtxB3cCoWyf6m4dpAhGIUIqkzH3euflJuM9r7nLTzBlEzW3s
KPhXZWYe22rM65n7w9lo9p1pqOWJrltlTz9EJH5o6bEm3BLfupgh/3yWLdbByUkQ
22eA3c/Ne+d8/dZBof217MJg/zKuFUn+CLhr7hZjRFQySrKRGpWb85JPtnW1ftCP
aCKbHqSJOc6eYbjZ/9UHL36cxCyncKQEkbPpp9iFQUWqifNaEViIfLvqUroZ5KEK
tfQMzgEUW8X9Tzb/trBP0wfx0XMTckHvQnVk/02OI8b1weSjV95cmdnc77zio/NT
T/CzXS+eUj4UPM10qe4ruKvZ/DMDVducKzA273jIixZ4PgLvtAEB7r8xRn57wrXf
dwWHW+F32Y8800/hSlfAk3PqKUMVC9Y6y3HOtOoDhdAESjwzh64NsEXTXcr8UWmc
hhcEBv5B5Pvv0P+3xX8j3wrLeGTso91lS3lj4gftp1IOvmZAzCBenGlz/QsJOmQ0
wB2IkO0+6ARclPJmA3xU7EpDweW9LTU+FDNfpW3MzGIdOpfcSnlxat+8KrAz5PHU
HscOR+op/ichnEaBGbMnqIjkeBe0ziuSmyTTWmf6KrXAp+q7wpHd9a+lVwnkrAOo
viQiQvxVu+Woy7VkJe5vyQ5anpVDz6rKhbVQXT0GphOecBK0WSSjtVhlU91Up9AC
f967xQNCRJHYj0owL3+qCptXrq8/DEHbLYFGNxG/IYiY99Eq7AqRc8einH8bXq7E
jlf2wv1iUFKitVaPOTR0b+3YAyEN7zxaiSIpLerZ+yigAo8kgC05qU1/3PUhQf38
s1ouvxv1JuR2efNYf3ce+g02kkRBblsXkEXe5NvCD8prQR+gXyBkem9M/sSXmma0
NBbAr6Ru8L1Q5vPP/pIsaNrLQM3CcPney9i5OVHi2oYVFsnHg8JiT4hGMlv9FewE
A4E+DFy2gExC/PvMi0c2By1d2QyC4RvnUe+0g02UQhnKOvluFrlCmQS6kN0A1unS
ZPdPwqbyotof8fpoeAC+ri2+Wklv9rJaESmLvlvR6kJOypPNvpReMoHevhJkjqbX
DSWpYv1BPjiq0vVDwmJ0NaWuh6M8YTd6FctXoSsaf28rR5EIdJWyOHnVVOl75dOc
JM1RlneFUKgS2wDI2FYSjFq7difQDVir5Wln7z6Jiwn1MdTslhvxEBtOlz5pklRa
dVPWKlgb6Tjy595rm6E2cvj2VParKKCC9ZuByj1yRdFAYBl/aMCbA9MIk5IKhAVM
Lk0LoRR01hIZbFoR0Gw5wuh5JeKXxy12CZIjteUJgiCn0/8SHgc1v6cK4KCUa3A1
7DkqksvP1xsjOFvNQ9/ubn/gjgvN0MVpHQnLP8ytexB0pasww1Zd6BuzFQXDYoWY
+Qyf0/0Ydb1jTXoH5haP+5DGmBkZje5TKqONOEwuaxiE2sP6xTUMgBB73KO0BYeD
Ymp083nv5RJLzAXjzfAkrYIEfRJT1mmpoRMyX6s2Z3NwaywoONfX8xTaTw5N5oeB
xABpYUj5gSxQmMbrdzaveUWsUBCHpB8EzJpPsBeOoUZvKp9ZRJFXsU7twe3uxJNv
7DRewuUV4tneRULroRb38555f5mtjoE/PRCLHqbsvJzDRv7MLB49SQXwPkheLxdX
b8c7OWP1Gjjev5AMk3YXIULe+tHISnYLgUvqjj02JXyh8dWlLZ2uv6e6gA9r2VEM
71vvE8HqPYpxWNxeXyG0ORSPjh/g3PMazOD/dpZXAdZajFfC0oo22ScOMwG14lnZ
wj36UpUqSo7WKnK9/4GC8OFs5gR4Mlpzi/97SWaF49ilPYK+5KKVw3LrnMRvVVeP
BrqGFuT7o+iB9KF/KwHdAWIF1SydOBR9OEoZWosx7IjvTDDoxACagbBUTIwg+/4V
MN8Ytar5+nPpOZXWfq7FVdzLMmF9QLGQs1TXYyp3NWBfrEAZxuxv7K4Uk0T+Bm7o
wLdllt0jV4Yb9fJQbtu4fWOuTUAqzn8TFFb/ous/Q9tKY0ymyceANjzwTcOTL78e
QXjiI6ZCKReA7JDziEw+JFv9SGEdH+O+KlIKkD8qP2IsNmNBjSHbBUgKMJ8SFkaa
sKjN07ia8TcqUt6jZ/1oQLFtn9IvJSsB/BaPey3P+Tx4Wh46pqVOlPwphi8bou5x
BTQ6y9xGdZEgSen1pucrp4W5wSZSpYDJa2ae+D6aSqGs0Kv/Pm0U/f4XZAZ4M1T/
M6KLtA2lakQsg3z7+Ijm5KJCmbjZEBnYmw9U/tvB37dBjBM5ueZea6Tswr31wcO+
4/pLTxOaneMnX+Ql6gZ2uWc4kpd8qO6erwlQs970OT7bmTAHc4jhdA1E3b3xBVRu
/YmXP7egQazkKvz+PE1z661IYbXnmcwNstABoNspth+NnAph2/So4K/JERpB0CZK
+nPfxNbssfR1fwGGMQjdjtwW5+AndTEXolvQQwpeBWeSh9XBQltu17/mytlQIBL4
UwHB+kXwyzK1AZxhPrCTYlaD/tQ20ssSEpta5x4DvYrua0b5o6t9xdnDKwM1zSt4
Ts1+gA1NCjNyKJ62yopW4aWGuqGa8q4uu3WFBhtatQUB8608sgQ0h6do2LPNUuPY
kpXX++t0mZbZZ5zMmTsdZbgbpaM9Kf+4riMG8+0iTaNvtxaxF/7W7llA8cbAkBST
iLOHJPAcJH9Vo0c37zPnucGmL++X9eI+mfpg62+j3SBiG0RqepLg0gldwvOiaQ4y
IByYWOY6jBtDU+SrJEJlX7mK61TC1jyH7exzzhROK8wmLlRXXHrspLWiSO1WIXmG
DflgYEqqGL/LQOJQXp9L29HSrJQ1lxQlgwd/+Mc6CzUbGve9JZe4f5XMV9UhhiR8
WRad005OlL6GXn0rebahe+OJv7lE2OMgVpg2Qdj22ixhcIX9K8/6Y/G2//6DZ52u
28mWv7B//UZ8Su744SPXJ1kA2b9XkRjQkSSC1vrdr8vRP++kftGVSC8Gd/CJlFvK
lI+TXLYt+fDTx3Db3U4cXyJ9mcze/P+UmsNPxCZ3UBNBV6qrX5uJM88uWiGvor2F
81qKmH5CF49gVayxOIzrdlGo8floG3f10EZ4SA6xo+kvwOpirThUvBo7dGrQDQrO
+2vZy8m+sAI/Dg+gOw9AYmAazqw0b5Y5qPSx934S5YFvfO69s3UpEJjtAq1hQMKR
vEDdtkX4QaDDhPRCEGA+DuAXzZ9HJdQSw2ilvUhSR850UqE0m6H8nz7jOOnIH8Kb
ex5mXCU/UtbjIV+mL1i8Zl8w5IPeagzdaTspgQM1eGHRNJGtaMskvJePeXe+5Jjn
yCGG9zc0dIHQOWHWGyUjOZSsAV7Q2rBNCJRVFNHxRS3E8dwfcqrrHPoHv2MUMXlY
Aa/2AuUtzu+b4eIflzoFfzK8rAHZIDkHKgNfVECEHc/f0aMOM0NLVqm0jxZeLWcl
pieUEo21/K5A6lSsgu3YeB+DQZ0sDJvt3kVDGwnRELUNDRS82gycS4L8sgcqyYfp
VtvBgt0mDWi/M742xMaXm9fWEd0W6wdTcMIizf5YO+Gqh9wF9hvfWERtqPdn6rcL
rvJhDlxCK40tUnTUaheQvCZ3QExPQM9N0gZUQcIy8NRtXzZPK5Fe0t53xbv//jlW
ZIxzTXcFkA9ZwiMhPjVST/agceFVq+QolknAh2BKI2tiSriJgCunh2AkwiLzZ/0D
j/F0zi9+g208d2IhQWJfR0laSBXYqCcin6FJIp17gT79R+keKgp5lJ2GOBuHkwhb
jALkfJnEypjRyzlGKmI/icID2vxznmQe7caQrFCze9NooobJm20cRmGKyXrGwcHO
mdU1pEx6sVPpQGP3wqMGnE5n2VonpPg0JunCdRGuO7ewAqNCQQTGfeP6u5mfQOyD
w24qObGE/DcVxnNkjRHCDnQjbrchYpwgTBRTOdwKkSNAJqUrPVkF4dSMGk+t7ww1
G6AdkhadTUfeucQmeil7DVuomPmPutW2GQsGkaO8zMrU0RXjQIjW+Q5wizJhqvJD
m3tG1gBNGBsNUvg8Ua9piFsr2rJnRFefKctVZee9hl5RPlm326ffZnrh0SZqcUbL
q/P1NwYhlliYXlt4QZGwp+3l1hlGpv0+7NH40mk162w4kHv1gw9jda/564zzpgzb
1zlnMU1I5KZt85t6VUnnERhix70xMeYZ3oNLpN7w8IGywhjS7+NkamiPX/VwyyVI
0KjVUMCUZKsY1yyBWU/7LokN1ciMtuNT1kU9sqtFlupbJimzroXHLfZ8W9yzSgbh
I1wy263znURQAckzOeMIIyVh0gonoCQ1TZJZzLmzzvuecdKOxuUYL+8787mG3X8s
f7IpoYQvZuWf7dscHWcM8RVDg1BiDtlRvLNbrSiMJXS8cKvtcbCH0Lj3mY6QjVUO
BsT+QB9o4tz8i5R0wFYZNdfJSAti4gk0UAlXDtbVAelDt566k5TtWMtuA1DqpP2L
LtQZjssPcd4V1RFRDAGtUrnlautPyFReOq847bGJH+iQjK7rjeYOHRmgeAvlLTV8
iXzJEx/FhqujGAWCOfmVq9I8Zhgk6wAd+YQYf5CdY9wRBH+uaio9hvkRpTzTq+vU
t0UxgvoxiMUeEJHbfzxvQCi+It069BAOG+mrDwYumst6xvmbSHoA4iqRcktDdTeB
9bIXI5dXYS+h7/LidCe5hTYXojQ0hyX9VNwrjpW6rT84IJMIGnOXlbyQiYIcTJk4
ELeoG/tLrHwEfOcoPkCjR/qgNfUVdQtl7q6rETN2mIdYUEfxh4590xu/HDVmLrLK
JQwkd0t/MyKL9hX0T/14HzXSt8agFrEV55JkfMOPJyXmdQDx3ZCIcw+eEH8pD5RI
f1FqIZmowND9wJhMDxYQ8L11LZ56jd872kXxbGwGegMnpvh7z/x9iixgsyiU+Thn
ql4qagGmvsRX9lCDvFWSQ3+fF18UvwzfERknohoB9oyo/LuuwGSE2deEM27ppiRz
8Qslnohv7StmbxEg6L7iCD0kiHOByvYhZ/n0glqVYCElUgmX6A0xmGO+MiOLKhS8
JZP68l9wOxgtkMy31vSgrWDCvkeGWZN6/vi2UL5GTxfAW6Zi/Bqf7unjZj0BSy3a
saJOWTg2DpTfXh1RcdDDqpAfaweY+l8r2+OvSITcphIAqNZvkRTLjlDUyiLguyKl
LPc2TF15rRwmk6Dg1CIb03TstzfgNWkoMtdV8Z37IBqf5as07J8yOSiHNm6zg/p9
84Ikk2V4sPfb1Xb7h5cl0SqGG1wvR0CYIY5EUg2qk0iJksBTEn4S10sxeKeUennZ
wa+vlfZCckz1jkev1+7B3jE+HpNmMoD+qam1KkXIniZpcSbWBfsrsROsqnRtDtHy
dyW1LdXOxMj+Iqd/u8QL/1nwoftycUbLintmE5/yOoi4HtG6Ey1J7m8W5R8I/GfX
YoshcoixnH9/5Z5koKKJAMmC7EnVAa/QrGCJO08zuEjqtIKDwQcjcMhOvQLy32VZ
09+WQGwsNW+zN/K107qBkWIGkdLjzWlAaH2xyCqVrrfg5n0ejoy+dSkZ2ElBcoqi
OVK3ekFLwDkAhF4WWVnognhXzPEVi0upqS0ly02j+GvcDDm8Evg0K+f+ueOX+JRn
tDEv523UtCENT8Wuf0yfxJIipPVVEitn6hGJyY3YDhxCK/xc+PM83RTVTuhc8DjE
JELHGfOgo4nsmpbwKtJ2qA==
`pragma protect end_protected
