// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:36:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VcuJLqqRkaZP5VjGxFSng0K2mCRsNEy54ZU2y5IThuiumBxnaQA3eP4Ig9vsKC9v
XGinJjgfAdWUf9MjTNqsUca+TQwuu9HNK6IPrpXGQmE6CX/2Krk1WN5PQHQtb/vy
OtQbU5WLT9KTbFWkZR0JAl20yJmsF2h3A/Vy+TTXjRw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3584)
Sh5m7l9SaE7i3yZYWSZ9h9Pb/GRicu24Io0lvZhlW/Z2hiOjzbXTwovjVO2ow1yF
+0tBVD3gfmsarNoJbhSqX1Zbjyo81l7zNKN0fm4IEGBZDzCOPtDXjUToDSU9DoMu
dx2D72RUC1vMP0F4MVDX0ZCUzguyxCcxE7kp7YbqG/rnuz/UrT9dOYyfogxca9Of
mrh78qZ4hdrlMntkR1MdZ6zb5vIzNLZKcVSm+4MUiwHlDvipHmpidzjX+XiiH9QZ
lqpInOEAVovsW8qYQG4gPI0K4a2STGoDxYmmliZu3LJD0Oh5bzMtzux+rmcpwS4j
ATWbuad099KxX9Vn0LGdYgoLkRNorPz+ffXZGfJvzTT9pQfxDNcbkbZ8rOUaGx3l
/Cd3OuVrW/lpvPfmqb+eNV7bxTDUdX5EV91uU4IIRTvG/LNYJpWHR8SJeT+gBrNO
3bg01BusvUflpt5zIguhsWSzfElwlovITrX1MZ25XaG4n0ZNP7LbFuc55xEyhCUC
1cKGj6XFIBSMxBmYAn1xocOHGfs9Q1jRJmKRABJWAXgpbpaccHhfVMLpPLu4M4LJ
u/WaW1QCq9JoqgMi/JA+l8EHIyrMjrcSATwFrVyD29uS+PLYSwy4TnIphSgP0c5z
E50KrCulgp7jd7thq+PFavNVR0/kIpNZ8WISHhk43b5Cb4+qK+pptccBKOpUQWNZ
wu6qssbAw6iKZRKs8izFhvfW9GJUSczyMQt8jZY0F2JdZ1JEzHW4JiwL35mqNHHx
LaZ4W7hz+FNILWAQb+1K33AqkLjY95c+y+HpEqJ5U+0J9K/BZvuz4LMd1FQfzPBO
HCu3TVNNW65f1wvVngb7H3aNzXj6npUFtcx5WcStcGxfS+SYYhCls5WMI/CNe219
LZgAAu1CQQyJwoNCiO8/54xQRVKLS/WWvL0YXbgceWUreXMDpA9cy+Wnyu8Thzfp
B5oyg+EKxGreIu4wSDAE5ElmAXY0oBwMCEupLYLB4jvcM1sdNQxmaT76NnpULiXN
omGXubcetlw6ruU9P9NNCgVQHrIHFniSNv4K/oAqd5uB59svHB0FMrtCF/oj6yyF
/8roNtKN7JTqtm9S1nn7WvHI87rlGbYIKuC4XJi8fOc3HHLx/qYd1D7J8sGziwnZ
C1lyieecJBeI+kogvCjuKkDIcwvp5zyWV3n/7zy8MQLwfMNpHMereylnj4hKGn3m
95LyIyUDLfeWyZ9bOEOYNBu4/xVl3bNxm/alLr5sLFDL4b06/FG/wSSTFoJK+9Na
4Q85Kys4gj/YfztJXub77PDXzKPMe/XLDwASrFr40TQNNLThY7IhfThTImpbwELL
zl/anzu3zEt5GCq1fJBNQvG+FJWixUUgvQC4TilpfgUn2tH5PAy65hR9WTer4HQv
+OOYUlMrI+cQs6NHadpXJyr7z+CjKVjacR5kbjpnKklKORMgBun7qyfQbS3Se2yH
ntaEkBYH4XLYQGgTzDzMN1skhcjteHbINX7lA6IzJh4zD5YqFp3/HALYSOt9i+52
R4+X3sdODIXAtc7wBfrv8R8HamWXXJHutQNueGH9IW6QxfvMW+OoVHufpHWg0EWQ
Y4iiBWvwJ7O/0S+GoDE+l2Whf1tfYKBHXtXYgbraYNPeRtosixQIUfvJPU/MxsRI
slz5diD96dPxV39WPuqKb9oPEQ4VtRmNYrj3xPF6MSihBtJoxe1hbOUTBVyhTnB5
5dx9rj4yRCSCv36Q16/ySUp5pLhAtqjP06co0qnkJBC1bMdHdV8U4d9T3Xl6ikjG
N+21bnRXVHym4noWYZdJ9U+dGxzl8Vm1Wth5Nki5ZMotSdRFZaJ6rGhuy+Cybt+g
msWEKiiCwN07+5Srh7xeISld8JykwmWiyktfrOJH6apE5posXS2pyjGDXUznj3gY
wg7ExJu53E8Xe5jeFwYcV+SJQ0EMarVfPTqNg4uFsAQed4VS36dJPObr1TYegVEH
ukXEjr1f0gAGtRQ7mpwn/Mpe8byRQu3NPJm1mrh5/QPmsp8JJNSzsixZlpPFCNB/
OhsNpAXyb7/ojTOeglVGKLIykacpcUlaNcqV4kAalJyA5jRq26jamhtyIoWAfl+A
vImV2Rtz9rmIRvLkxx2QRjt7bj/Bkc8IoOVtpdkIsdUotYeZzv8FpbmMvFYMjkut
QbSU3gi2jTEYOtAsSmuPlLgtyyX8n92nXCr99XALebTrR1UkMexDeAm0EDiVCfzD
mYGPVGduUFN+fLGkpggevOoM+d5I1IUdTs34u/4VWhi/fbP0vMi8NfbDtH4oasIC
iwF74X9SBwAn4Hv5AAqa5OJMtTZql6ywLo1Dcvzi2j+rL0WnnVdHtH7hvR+W9L2p
qMKdT0E6SXyWtYD24jUBVxfQ9XHIWtqu1D2fTAmA/k6aAbe6u9/FSMOOagXowpA0
sO1TscdWs25Rkye+eI1J/eSjXV5mbFYzBPROcjsw+4nRqPmgQOVW8vVDpCWxeNVS
BQA53wf8ffrfle7ij/W2bymZgO583X65IG7Fax+UvH8yzri2qummx8rQKAETp0Jt
K2oIU602Fd/EMWKjepw3qegAknT8z1TCVjcsj4YHs4GaCOlD9qHPZZYM2SP2Ca+Z
8Pt/gETy/KaUqdoM8uaJjuhT6HDkdMEEctAomdiApMeoYRWXul9jMBIyM1cDf6jD
zyqso9+xGvysVlpbWvpKBkMhkBIXHMtYmZzH2bqzlq1TGMjZDP7swICEKMrGcOab
Q4sEu9v6XR1qp/SH8bOePwLB28Z/YfCOUDsiQbX7JgGtLvKJmIb/IonhX/RuVgvg
ychU9kNcfjh/TgFm3bIERJ9iNOaA5AY7/LQqaMmfxbP+1LybO4VMnGM/SW60OkQO
GBbDC38gyvr7oBvlQ9X2kRCi2ylvpyfk3eOeV356Z4YygbNh7BTMXGklgTwNR0z8
LVZUli/USFlDfHR3qytBU2zo0aMasJlwCMf0jDTP4jsBbzXeMAY/UZTamQl9Y1Ui
zQb/eNqOXgytucC6p16TlRXLNYZfqVA+YVvRrp8+oep+nw+qfqp9u+LAwl+ujaTK
iF2hmYCBlKRRMHKtSuQaVgL2rt+vELimieGIngTpAkKvaADikc8JjKozY+EJbzgp
n8KyFQKyI6ixg/cMUt8HRg9B4ALDEaxR7TTq+oeovVMa9pW2dlVS43SfQ5wkFLL7
1V8AxGptSJ8AV4ShXd/ToEzEtQm6kdVpsAI94p6wmYLTbMqeOwStycGWFjkCm1ca
3HICg6wbSJYFtXMWQzz2Jz67g8Ugndm22yVRGWVzXiluBFZkjTYDoDGVX5fjADdW
KDi7oYrBrXPLNkwphEqxHL/92GywlDwoOEXIw5dxK1bP9YNirSBwQ6tXHbqRChId
tpD8/5DdgHK5NKbr06sjRDhGNQ63gqZVFU14kUIH4ikwH8/yIcJ/uiIiSiDTbJsE
IgQt1WNd7dzAS7V8NIdsgdGqP5Vgqfb8clwnvShOobPJRMh5AzACf6lx4a/wODk9
DW8recmLdKxx53CufxrBnmwqRsv+ZCUQeffhbvqwMIqKLddsBi1cFeMZTUZxe/Px
7UbK4Mc81bnjdf+ujB4H39JrcTObTixWE1pWunqoCkixaKNTHDcRCgCWvamS86VY
hlgwB7fN8LvBRMxC1xDe4q1S3gKd9rYmQej7DQu8eKjdLJr76Gxxe7w1dRq0CTyV
jaxkvv0KZrdPYErUEqWW/b1GBUiqmoVr7JkX3k03U6BrjGqU0JRPhoKniMFZqoTy
VYzGO6f5HMn0ainebtjMHZE+WmddXniOP7/R6Pj4DYS5f4IHwTo5tG/s+ApVeMK6
ssRFABHRMc7B6YFQD9IZAUtityh9tLNg8BH1Atuv1hy1CGMNZp5gYWhGj0xTPBD4
iZFDDWedfxbWDdTkWCn1tNgsmm7iii0Sw7QO6Jl5PaBvYKoQXigkgBQEIRz6x1l5
s+0jTV8Fn0Hz18H9pgB4robcEDcmnRtnXaMKSvmpObc3lHG+peSdJh2Tq3YfSefB
c74g0C+vL6wa9ZNbm/WYzZeb9pVvf5XTiSFeFjMwuDUMIK0IXN1tRMiaZKpR6Hxi
R3ns413un7OrGcEfoGnecBpi6TmORjg8dHTDC6RjjrZU/1VziFx74hmA3o64dqtI
H6bJDNqGZdDY1VnK/UazSa6btOa5Sv+n9U7Mgr1YFaoy1AEnaPruBaVJcVWHt9IP
fqIfjJ7wHJeBtq93UQ2FNzOiKnn1axpiicLFuPkEE7HvOoO3790WbD4vs2F8C5xa
CnVG2ADmUxS63urA2KfXE2Q52k2cfS8twukLyZe5CR1YA2l0BPkfYz8oZROTTMsu
TBEtINM7ciXMnqUalUbM/H603wPMPhmlgz5658WtleaQUcLTOqJTPDavv3XiR4HL
4uet6hEW9ouO5s1yDyksLLMA007YeypJu0srEct40s/vIyyJ/ijDkzWrgfdSO5un
BnblNaNG0WuaLK+VrYI/nTYHlCOYe3lYNuBycbybHEVss229Q/tE80WuwNmxNZuB
1kJ+HJ5IrO7SWLExg8oydwBohnBiDSNY4si444VCZo5TvOTe+tWiRz47DjCfwg/v
lz4tN7IlIWp3IVmV3vAHBEP370HhO+CcJfJ7bs1T7DfsgHlW0EKjDP7eEucJqf/M
k7RejQwlz1HGpls3DzOjbaH2RXnNueLMsPJLJ+C8kuXOTFfOvxCPMBv0/UNHmXRw
QYl8rjxUPZN5fNgkRYqMEV64oDiFw6Evb/bZMCaemSI=
`pragma protect end_protected
