// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XHQNX9/YaQxRTxPQydCvCpBmLp9I81fCWnFCKINbUO4GCCn10qERRb2BLlSS0YVF
8K9zLf/upVz0R5HfjUbQfxHhkLcGvQQ2AGt9Ob6Jt5bqn/68KwhPeyq/vtM2zPCO
q37Mt8kJqEDTNFlRxoLbD6cDlyEpJdOy403pXYXDEVU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
DJ+HdSWMiBy70Eg3HCDCxEH2a4kkoLzmZNT8Qqbh3ztdhR1nsrbKjzUZ6CDppij2
0BvJuttkL0qyKAgVbOkv+jV/IUxZ0wiUo6fe7j6bmbbRv8U5UusMUKsx2nh7cPbo
4RuGVgBMtPURWNCoz+HQRAH2smVwmdnGx6yiujL65qszbQ6AKrh/5tk54hZKpPEk
SZ+vkqNsCayHYfk8SVot3R+OVf0vNdURcjyv62OKutWL3Moc5FbynX+ZRL1LfkDj
8pXTfvRsPHcEAiioInCldLxJiNLxk9dg4lA12nGOYekep/HMd9MafNZRAWHQ+mtl
k5yGVWjjtt8cneLX52ezTz7ZWYL2jHVocAL2UnFUQRfBec7yPy5/0+V+uDXvI637
CZ/vOKdA36IntruGAUfcYFfVw+68+URKuAJ7umt1tIQnX9ZYf55DSd8Ma5hvON9J
rSQ02xKZHbCT8JnA76AFX98Za4X7lPY//wrycwWSPPwGPYQmBx74RQvxiu4lJfEx
neqbw9Quao4TPwSfaAzYrwc6Opy7yAgPrrgl4QrXVmJsYNlzfnU0I3PD7fZRju4f
MgqKyOyYE6mJKTJyb6IzQ4977BIGlptnNn1JEvqP3gRoHDzykLKwEQ1bBbW6Wqqv
p1WcGARXNa5IjKc3MiIKNWQ+WBwHdZxmlF4x2wxNnThCsh/0QtuXRF/G36rG4s+c
3BHSm0JbBz3//FKdhi7eM3T6R7zyw0dE7d401Wb4xnE+rBPM5GhJ/enMvUFNmE7L
KOaHZEHJ1BK1iULqx9idjzfj8Skw3dm5Oc/jpbzR4BonsSxDiH7sPLxYQfEIFAXF
BpLV4jyv/HDvf99IybNsdY0jsR7sL2vhlRfsxyVHZWsgirQcQgddVSeYCzzLlkI+
K1GU/iB/UvZ0QOAZfPxdAMrX1TRwM+p0HhJiHvMBMBQfmQfCgG6flYcvVvL+d+ax
GljivaBxekXLf3CUO9R3I7GCbc/yZoy3yHi9ek1oavorR361LXdJ/g4tYbjFMlBn
NqPgckgqmDEKDr7497xtwVmm1nu7sjd4a28iDk+6VEjslX35dP4I+cWpdlK32+Q/
Z+Hb2hWP1rpoAhN2Eaia/CwbdujzYKjTfxw3Ex1l9muD3iCHegsS61Hml5SqasGK
3pbg34N0kp6VO6Od3iDzCsFB5M9Cuou/t+6TuRKCVEKmKpcXuJKJ/36RdEzS+yMp
t4bl6ctWQn5I5KYNI8cU7wtx6PibrwbLomI1/oRcQGirQe3JQb1T4IaLE6i6hlRr
rpvLII4i26L38GLks+Z5vl8ExQCA0QsYNrVAJylgda5a4gXuDhaX7Q/wKmnkZL7t
CzcNqrHTdWkooV0JVklfbzWX1m5Z6MtDBSyGiEueYr2U1cSTsilVCg3rN2cxWIjn
f8Y0UGwPNllF5JI+ortwSxv263paWc+WWVYlbDO6MgEt/jtu+hCFRNLoax0IF0wb
EOJAKGvV/Y2aBjw9LpIepTQiRG388I5Qq4V0X/MabLJpwkQvRgwc0qiyfieLApmK
WGZRusypGIToGJ9F+NRIGQr3YDn1uCZEgvMneRlBOf0ojkw+OM2m1B21QkhUoSHN
PaVRUxp5h98podBkVA8LssuuVzb8NgffjUlL5LkIwW1Q3w7UI1OeCL/PzMP+KLXa
1OwwrJT36WS1d+8zRDSZeNk0jgAxY+DxcEllFWs/FzeaBV49FwyO0OIrc/8bfGi/
PQ1o4cfqi5s7oh9VN2E/GcsLr87OVNX6RuaBzC5/EP7vAwyJLlNh+cdal5MKsgF4
tHQc9Se8BOQoRwYGczA/6lstPs8DtAGp1Hj3mSG9QX/ivuPogpVWn+nF0oVYAQp7
1ZF/KL173ftB8326BFvmiXe6AHSWlW9znPa+91WvrGkntG+p1TPyGXSbTaS3s4uD
uu3TcjouRi2G4pEqGiGiCgVnmx1AJ4BRMU1cm4kf5CSfbROZoBR3Oo5k83mGi866
M2z4WLBeisRAP9piGx5uMCTiQ9yKtcAC4evszinZJUzfi4YTmwRIbuQ2RLfXRhOM
i6SW6mgMtf1Z5aw+edjS//+jN6F6Ey1JEpI3jX0sRPa23tX/zGbO6fXpKgInRUSH
7Q7u5378ItFww2j6d5mxPxmis3KPMOWHfFuShbweQt2D9LcDrG1iqop0Cif4pJ+5
n9R9jG9C4P0Wm/hP4TjtNCvnswPxO1lkLdc7Hq6VTV9RXF44ednTMeYJ+uDiO4l2
QPO3Pt1PKob3wdnfWS67GpR0ERsusZV/NxCFObKaPMIGbA9NuMTRkdYfObokqIok
Fh9W9U/MP14pviSZ2h+OxhzBYZhI5vkIlNo2C/GrSScMX+33IQbTWDIVq0kHe4F3
i2LgCvIM/Q4s3nBeuuJX/+1Xeos++0s0PJJ8F0hn3kdviMTIHcW89dZXzWIHPkFd
LLqKfigPEcoQ0qnc6it6Wm/biPnGskRvICV7HNbkmLQQO7mlx8gnsP4eGovtFGir
ZdYq8uSnDnzxoxSKsNbh8cARzM+drbFNKi7z58nRn80Vu5ZIN+GX9psFhpHCOcqW
16/voHAN27dTtRhhN/0vXUKLxsM48W5WifJ4vN2giLhCoa9dwgpAczlunY2yACtP
aZWEEviJgViidyPxj8O43rW94iqlSlPcYzo8GDSVwMAyN/zcYXPlPTItB2ZqqPqe
7QtEruTmI6kLMmq7t9HBH0R5w9LkAVZRGFmgfXz2/JcXCRQT/C/KsVam9ry8u0FK
Zu2dwIDaC9WAKrLLl70dTJdwSP7/M9P8uHeBrPd7N0yCOY+VvNxTPb3sRTEWc3pa
aaXGjCkvB11ef9sBhrCA+RATlMaFjn2x3lOpHDaPuzvzrtWkJxWJlKYMCA4nqoeC
d8ye53KA5WeDSJy47SysbY87lLkxVBuXBPZtaB/gKYVZZLrLPitTPGnle+3F36Ke
3lhEl0bpe/ly6qYpP6Q3yNU+m8vVZ6CCEOCSH7xKB8U+MHPLe5oChtkMaW5XPMoC
w0m2byUAtPwoB1aOasQMUxaxA0qQmi1SGccWl4kjlR4MQ6X2WGweGCCnjyzNW4Yo
2ECA2g4r5E4GyqYrJoSyor3YidbQKvPXWa7KyLX93qKNujH6nUGCWld5f8Qt1h51
+hkPNvmPY+WSVga3oY/oyGqiUm8xGV2eDHOwdfLx0hELyZldcveiyMAVXMTf/Fr8
nUCvsvjN63CPImduObrjc99SOA+KJnx+ExziniFYuDipZZYsTnkY6OTL+l2Fpmr1
cMCJ2NYDS63cuqGZNuIh+JbUh/cEkFa/V3+eT5LfRaidRzJD0kIaoX4dlMV7o/ud
EwuapGFh6D3cVzPN+Ex6IXCK7QNV6DclQ0pQkHlJ7MzrHT1b3aFMxAtcznq7uWN9
pHYzabBaQznts/PWkihDUZB4RSSsweYpc3bvghxWg3Q/xrEOa71z+meYF9Hhhcla
R3BfR7mx0N44YqVAXwqXDVaWVO9SwO4cQ/m6tFv5nFn12oDlA70h9zLqocFOmcUp
60U9212hKhoh5+FQNJrXBrwc0l1//2YVo4kXMb+isUdsoOTUB/pPY8p+p0JJbFjA
WFUqtLStWZ7pTkLdiZ2VeP/UjHYBe2kBvMhdVsQweLEFFWgdsnlKY4Km5W5+g/vg
Fw1FYxlSXNHVPGplaZLV03jyY4Z3k4iFDFCRA2ndxmpsbDRkjdq8xNRHC7ltLceH
VdeC9dimZbZR3vhVmSer12tHdi51IcYZOWju+sXiPZ8oDpfvg9b8iJtaXUIbPgrN
j2r42ThRdZUDsjO8W9RreVRTSCB/wVWzOhe0MpEBQcY0QWSLPLUNQbuahnPTFypR
AnxwHYrqyWemGd36Jmpb9+BqgTW8HWtZbuhtfFcK6H5mSxR4+I3nubrMTm0dDH2I
z/vcMJzOwTMPNI7etfIGT8XtMUUa36Fux4WYSaXgP2nE3MRDzTYoTmokHBWKXrd+
hHNL8uo8NZy9/So+6q7SHxAjC7MHU/XBSKO4QEGtlLp8Ekdrvl6j92mQm7Ur5Ech
ZXocIH3GUsjS6pkipCkFfkkGEXDobca5EB1EclFGcjYfwtwnO4v0QYX/++quNE2o
1K2hme6Exsx6coVfHExH1vOGbkEbxwy54+3KC+iYVMYK9x4f4gHLuwBeRi1TLe7W
WwmVC/glGvOL+iMbJuBYjpHAtVJjk+0srqTVHHafaVhrALF6qfmMlFd/cBityTUK
8xbOD3vwYApNxYtIiDgAV2Yp0bsuato6N0VQ7dEFivThd194sfyMkch6b/G0ggPX
qgeLDw2088vSzFNn3yxJpKL2t+WxkC9D+4lF09p8ykSuxxpjyh+EfIp01Qwvvsqa
iF51+TGzNs9UeezbBxVaIJZESilu2qv58WN5ZNBKCQtsr0DO6SqpSGjDyk5dQ4Ud
tN9s292VURQHoVPq5qUF+oPXan9UvBogwf7Gsy768XSKwyCCvYASRulDdLeTIJJT
4isk6rjzm7+z7NsyYuV+fsq8NjH9B4YqFkfkAbPsHSclOck/tfFF18kxdysKMmyU
lg7JSCNintKAU4FNO9NFXxgkqha9mXTNzSVngvtUwctsEWEqZ97jbUwH3x7xZx/g
pC+zPvPagVxSmCrgMzMwvdNzxZhZWiD99UeLkBZnVcLGmmjmFUjIqf6icmAeBGyb
VEcvWQvtYT1go72YK74C+CujgdvJ1zpSWFN9rm9uznAsKpaYFtj2ddQWrzNquyof
CLyxsboGS46ZfjP7/O5ObRTRW6+MxgBy5/lfLTnYXcvZrfWu91uekWQa1LdKB93M
vbQNEHg01xer9/ZyrUODBnxsob4KZBN3miZctcbnOfSdMs1/xp9WYCAc4TzvQ2mk
h9NCPdyW4my4CAxRHvGbmAHmwgzw590/b0ameVn9Psiv4UeX9Hnd2FZi+oiZoavn
2VKvmPpiF+ZU13zeyJ3vdagXIkcDmWiJzglNx9ism0SQcyJ2mQoDsexBUEljUM08
05Kx7ZI+v58En+R88yvlETOYPnH0Z8JVH2GoXZDgaramrEw7ukjl4VfgLTQCIS3V
04aPfD9oeXS69JjnSepFduRNTVTgyxoMOwxmOaMLqHeYODTLTOZ3ttma+qZs5g+S
2l/jzpKyRFQfUTpDvdjOdOlI0vkmzuOcfQYnsXpVFgM6bdhUxluyYwV64qA2GEY3
XD1OvmbTcaeXreZTxTF57O8vAKSdf1wmzFM+VbdCPrWF0ESFXJ8YaK7riiDR9+4P
AV8na8CT5GktMrdK7w7SgrsVLVhLrCRkCxwsqRREbdxymNawcrYZLSc9toDz7iFO
xU/+Vjl0cz/i/ybGN+eSE1DB78TFkBw2y+6znJ+CJ+M1r86SUEuKDsjJsmAGRJ4R
7g77cmVSbQv5nkFnFpU+YpqDYlqTj99D/qTQCHkAms6ytJ4hNxZZJL2DTf9PL06L
hSi7y1CviK7NGdtwzj7anrXgJS2Ln/tD+nVd5GLKCNEB0w+0b4tn2k7gp/rdonOn
yKMYkdB98pU2NmOmnsEzkfG2ULmVfDyH/MvpSmJ8ffs7crtk++Rd6aPUFrkgd7i/
pmwU5GjWL8yXi2mbf9K5Iqy8fIv2uVlUXqhCyQtQ1m4y57IolNqecSEYi947n/9u
7BqlBiFaPO5y3dNU4ui1kz7o8aHOVXR8QwCcvVQFghUgt1uQuhUeEH92EWgICUQm
cvG2o75zEWmu4h2cCozIpjwGoLpIJPNkTzLXfKDRXk9lPjTqvNSkerFsXkw62AGO
qsGFY91kkjuCV98Vh3qIMhmdCUAPQy/HECAtJ/MN5CA8NFxK+yqAYvLNuC7AaOKI
+EbrF/0MaWsruma8VmGMNt0baI8+xGwAluOBAIxvyLdBRhXeSQ+0skbMJi1Cs5fw
qXmuZlsnjzxz4DAgguTGu3VEj/QMlUSbsGZIeCIvtl2llVBB+My78ZQPutygRlxm
zSmYXb00ZBXWMa7P9vBP77Jed9RqiIzWYchHLPR1xwZRjRvzdD+MHjJBXZ+jSiRv
BPhtul9T0FOdCS+1B7IDhycScLsuh0ov2ST9gSkXPckKxmsu5eJRdBpu+oYYmBxq
gy68rnr1gVq2to3rDj1rLV2m4XzpnCGbVeQeT/mvoEjmSMsT7Z/RqDB2Mtb1PqC/
nIbfqjdfz1N5LarnL5qLg2l2MY6nC9O+yjC7tjVkYhFSkm21DiEOPNf1JuWGZJNk
6spJvG9sCspQXaWvHARxmS6pQc5blCvgzoqMHBx0BtcGiBEUMONXMvcm/Iv0+ku1
oufrTyjARY6YQltyYVdBbxkplvfBFc/e/07XwjkwDQTlARyZsShCstd+gBrmr/fz
//hs/Mao0CABTNQqdu1uj0ayEmEJPsFczSwXugFRHXyZP8UoLByToEC52mJTQbUU
UkhKv2pe7kzAmttTjuh9lV419qn/sxL4HPdyvy+VffENb2jT/8ZT9gIkqx7CENeS
9pYbKhCYup56z8rDLbNt/n15GUBFKdtCwMOq7cLwVExJNNh1rQtbFn1nTIB8NNh9
TNwDGS3CFRsTtV/BkDwRCfNKGgAo9OM3olH7jfjSguOD/OMRTWMIZ8gmHXGyCwoN
o8w+L2M9f0qrbULHIh4gGnQr9F57LC6JSFIwYmOx2dXTSAUvHFHfWyU16KpxZ9kQ
HSmGkMo7GzD0MZUOo4jCFB+zuoVK/bkEPzhGPer5eAEZZLu6n7+Ve44xiP6kDftC
+wEOyp0lNQ+NnhKKCSiDh7E2ie4jb8ZUiTMm6nu6ItS9Xx8HG4zM6szidiMxyjxM
dlFsx5/t1hzUWO9MlIsVEiHBtp2NfcnFbyj1khj98AaSiBksF8NnBKri7Topn4ma
Y+kTnd/6UIosyNP7VlUX79PwYDNhk976KTs8eLBzqn0QTI1kgOEzI1yRSoDhRffn
Uy5cBDHEcTd3POZP4ndjyZwh2qR3wY/D4SZW6adL2K+rV7tas21aPR282B+yES+1
OmJYIhXzIUZaomoiiBmCyqK012MKqbVx/3omrhkdInUc2tHdZrtIkl9bx6GYU1Fs
Kd86EoU/Fj2ERqi8vNTrHHOtBAmXmVBuKCK6iNhwF2Suu3hjvWI7hObvJ/Qi2u0i
OG27wutYe0iBdRvgcTT1n+C2yBKZmCHKF62mIrcYMkrZRVdIgGyL3DFhfQy5Rzl7
tdF56CzUapub3PiAUf2Lyqv4TlAp7XBsGKALs5cionWcYTH3Dow+U2slXA5LKnnS
tnJqK9mUJ/iSFYdgSdW+B60bfmpZ8bliua0C9JW2vIh5srb9TTQUy5b5c9KKZag7
XYWuPVjxyoC74b+VRlRqaylOEOFAK/9zvAZ4rux1++/GsqYudODsG1bBEq5DUFUJ
Jkq00QOfh5O45oZ/Zu+EcIhTiX1t1ZHW4+xhXtzwbSVvFdbm6IolPKeFM01r1tOY
t5w3q370rp83KeuQFQCxKLwTUPwlhpUyKAZMMGB483nFLhyhPp6e2Z/PBtITi23n
Wm2vPwQj3MQJrmzdwzOM3uDbbtvPGxYo3rIY/g7xsVr2J1I9/2rWqCyzzBgGS2I+
h8Nfhv+f2ywSP9ELvufYItW+c5DOMHS1g5XJMGrbj07NDcsx9ILMvyAmf/iOKHlC
7WolBfdxtlgnEavifMjNOxMFhAZ9CmrHi6yreFdJ4V//OeOiHEu7WO6PtGvk568W
wLdYYlmjcA9aZeuvhOzLm1lZ0d0e+4y355xzqsP/S1+5PuQDmRSmmvlwimdRYVze
a+vZac21XAi0vyNfE6AChWx724beo73oiaRj8i4oTMZ2jaAAdaZ6rGaQzRidxLf8
m8asmpT5EOh/X/fgud4Zrjy1aT3WuhqYAMdQwFFyYchcBRZaZk46roo2PDJfusBF
VkwFthdaY5YoNpOj8YeuVMBOtaU9krlJ/tGr0qwtjnAxnvMY7QBD570zXNJDiRlN
PzlZCaa2JaQQK320eL7WWPPjQ0rJHWh4uSEKMgirAFsBjYXJrYYOQJt1l0Nr4eTS
DKMD8TG00R6y8UWlD/w9CpmyTHdXY1n7whUOf8cwRhfENQnOEXqmmVtuuF6N3Qx4
KRpp0B4YP+QkkSUBXnU0IBZZm22D3G3EP/EItWLcJMKmietFpPr2lnvIm/ap8/EE
ysxpmg+kG8t1Q3cHfHWOF7VxSGziesAuCUXSfDI/VEfJfmWFCcLGsbCTYnFS8H60
lcO8n+x9W1WlCZINLFk8wHfGaasuD5CkWaApu6bwjuSuK+7n0O4F7aYLWHlVpmHH
lOPr4EawaNhtlwMwfHsrx835A7FDRz1/O1DdSWHcshatIFMdZtd57rk1dxcz8SMc
VjnzGJ0tWTcPWrIDs41WrsgSE0dAihQYOL7oE4t31UYLDOSamj74i8KacAQRJ/Bc
CBU6RyR0bdHlkmgHdmbcgumanM9tF1PPB47Pa7bda4dQMGa11ksYv5+F794GSSH3
5uauza20I4zDZ/rLvGsbR9HJhWfZtk2TJOHP7HI/pG5r0VUixt3TmF7RCxTEtc/v
dC37ru1EkIjs3XGHQrQFtMi3hL1crfZS5VaEgcbufKlPypl19fnBoHL6paHtDOjP
h1PTRLTcBEFh8ZmW3LuGMv95yV8kZqlcwnD8Ugfwjx3iokmO+mDlhqslW9tKw7SK
OFcnLTbXW0f7i3/Da1PhVfF/FlSCY/MTPzXqn8TGa3m40KjOKoRpFM4JaEihixg5
CFm/uOdoqJTbMl8Yp45dhfzsN0Zi9WctbSgQGoEpOYpd2N29e3Ox19zMXK+Gogdr
N+tcBBcSCU7awe796UDoB/1xQzVXsEXlzqp8o10ZQP1mLbjeuqriPSTeq4j2tZRI
jnNqszUXVIPxm/Bw8jyc/KJpuHYj4HSsACmkXePJmAXFxlQpi7XhG+YdX9On1XJ3
5lkj3t17fXWSITgvKpaPtlzsBp8v1+K8KChu8sZ1mZwkLpMtVqdh83rfVgP5UA7v
sunm9BXgjXSnjPJu2Y9gL3a+cugdkDVEG1o7agR14wG2nFIc75WqnMxYBNHZLZqd
zFbNGc/D/kYh09/nq8lVou4uYnaSuFCRbRm+AMjGZlT1YuFLFSYC8UwQWLUZRotQ
VqVzW5+EaIavVzx78t/LAXP7B/hH276QtCBREL10rljX8+nFMoKmCWhBLQy0SlSH
bl69UDs41jhKREfdAmmok8Um8UaopwVrZSYHG1SvsaAC9wUcbFbasww2s0XKKs1e
ZprCRsisRzPX//njkeK5YWiYXNBzMk3J4FbZ8T5qvbN7mYOpsgGGtiQ7GSaf3APh
bJbYb/US/59WfQirsaarxsp8jy9hHgTyMvv0Mkjb2NZvsX8u6JmO5q1u4YbkCtNq
OeSy/zlEg9xN18Ij50ZfRz9CdZCSOOMsIVS7S6l5uPFvERTGxfxBbA28gXzeyTko
39KZy4H3VOGDA1G8qTCFX1/J8cJ7BM2bqqWAGTYCnT0peiwuzSYl9l6TkzfZJHCN
YdkXdU3WZeeBl4U/UpmqYhirgqvgIa5lw3euIP2bBt+WpIOlm3ExnosEZYJb6YzY
55SrdrdXY8yWLunOuvIhY2mmvvAKViL+gDuacbgC5u8ElZT8WZU4Qk0HYK9rhwhC
uQk+g7NYY8rKvruTJk7M+R+E4Z1606GvcP+WekOwV3NQH5h9a0WxTjVnRjcsjD3H
zLg/tmOz2HIXDyTY1qBwiCNmpm2LiP/YNXzUajeZsomHtfFjMwH/wuzxfo4+YBvD
86ty+f34si03wL+f39CBZehPXvPDLh7Hp4jlbbIH5efjg28inF4OA2VctR7CFJxS
G5NnSyA0SLGH0hxyINh/9czfMrijBXV2ViF6wO6dfPLjl8AlE7b56uB1wZeoLJrc
F/fFvwobd++f0RzoKERi+wS5zslT+l+NkhRRLqpE/AijMS5McHlQwWEzz1sLlChW
eIzMLgJ1Vd9Cys3WRonGUbA/d71AYv+/dHbeD68gUMHnUxyf8+wFfqyUhrsENwoT
VZq5PIUFr9Tsl8X/dqAZOBLRFCw5ysrzAWiAetfo5UurPlBPjue9Q1z1dujmtGR+
rMfyzPEGu1vA0iTniqU7e7hMJXOzHTYA+G3A2+of3IOuPduB2Ot6rBNU4soZEE/G
7VOj/AGS0tTtgq6jyzHd5ebI5dTYAY8es1uRoyUJgr7mAXvEyQd0s9iBpIFl/n4F
EL9EquQwDtIWfQDvrApRsE+Ahu7B/yNky2GCFyJXt+KKi4K4hqDIDsOSTQLWsMd4
cpmnMVwfVnyuXE9qrujFir8Sz8BM5UFfZKeukdZ6WEmyfnOu5opDKsczT/2vXCZ2
wCncGXdoi7cxIeYBLIZo7KLa7yOfoDeGzUsiCbsuHcbbxOg7Zr8CrbVX5fkKLFyM
jo522WVlmeAUjkpoOLgr09w9izxOyTm1At3rAdovJyJeJFbdNDi5uWPudBrPQeMU
mBrOPakjEDiJMKLuNA+iizu21Es3V+HqzOA+YQuWetr/cxcHiJw6h3irtYI9L6lb
mH9UjPgJPFcbhOhxCdP9k9z4gyM8+3u0gcns8oN2bvMdPHFVAFybcR6C/sp+F5k6
JCRLn8VXp6suEshYvWfSGk+EIWxSnmOPQkaUVsJPa3FNNdGReIiSljwGvtfoz9wK
n+S5w+2hqQcAB8mVb8/NcvCi2EIJxamh09LAGY0zoVjIM2r6TLlKcsID5jpIhT1h
R2N43KoH6No/BF7IGKds8IYjoO8/XZihpYcxwQ5C13l70VP/jpqYb+Nj/6KJEk3X
OrMBQTwxjKA+omVkH11XPWb4QBd2gqSBtuX8ettrj4KmD2lTHp/YzHUh+RpN74I0
cBZL8yvMLcXHA+zLJalfb4OGj6LYL1hTqN+UKRIvQE+WKdPkZ8KYi9kL0TZrP+G8
4Y+bEDVUS7vXPGBsIMkmsUSHD/6SFLdDr5dYx3YrImRXHJMTbOCcMZLep1AUQ9Mu
ZjJk7bTapI4Pj3twOvtnPEEM493lq/rW4I5IzP1eHeeMcMQ+joqhN7t1AyJ9UUdr
auYUJ+nScYbnyLRuTg+mcnIWBhgV3cm721cuI3eZnlv7gGg1sDCXhgQi7LuQaa2u
r4vi3XaxgTvcfbpKJMedj0mBo0sZqcLz3IN4PMtpJq0w8xwDkM+OSucDrwXtKEQ+
9XwzEbIWQqi4cDWYL4qfb7CruhF40DLskP3do1w7KG/OBMAgm4MTwnmyNyN/e9WE
R0sPfbHHWvynAoWPOebrCt1l1qFwYaWV9cdA4ErlCXrCiyG9nTBa20wxC5sUqP5o
sYsEImDO+m1yBL3KURp+SVx2czrlx4g+DSkYXDCphSc4VpVOg92AzNuID3w6Gnqu
pRi9Bld1q2xb7LU2EljfIcnBxVctlkpiPX3GMoM7i5Y9kk4ZdfPaj2xcCYLLug9s
lB3IVuets8vw9BLI7YcDonyjMDl+mQjvU4c45HxweLUSjh5LuatUg366MmtCADrq
UxU6G4+TpPSG09HejUS7S+LjduAEShArrHYFe2qSjIiMQpBhXCqmjfz0S6cbe4Dd
TV27z7gSuJdDNSFwmg+fkecXmjUMz0gMl/UKfT+Yo7m88oxbGF1lOSwrZVo1NNKL
VZ/HjnAQyixwtzImN/n+rPqOTWyPw9vQXk0qH6f2h4nTJV8w3nSmtl1NZICQvTm2
tGmlMg1GLz59Uw2ZRNMsfkdZylGwYQ/yimme0v3jA1vvESO7FZNB9helFK8iFLVy
fiIXYWDnatOyFJHVan7fbqTvZpDL9s3ljAFq5fgz/Ui0pXZK/geAWepf8cAdGwGz
66s6oeLMgrBL2NNQNIrlnUv9ybjMm+BewQjoiHRtKueNMgQu/UDmhngvzUfkShso
vT7S/g6NhIJBqWPz7flaqGKQkfUGvPMbk/iWMnRswOjZDQEaonZjqPSQnXq84Ly0
qNGdog2yFKSHSnVJ2f9oLjEeBHW2u/jyIVDG45ufcexGDoYhgzJiWxX4nDAkoGPJ
UJ8Fb1jau4Smh1sLeTuhrreNbCLnAGRVTg5ymEh8wIlG9+4s3XWCsxG7ouZm90b7
R7e6J9BtjIkgUH5Ori2IOGU/byQtwvR7ZAcCIkLIAvrW20FbmAA1sFeFefDGh/FC
zUGBdxXEUdQOkMyqJXpnflSy3VemVgpDSN1U23c+7MncxlC4CJEw+/85LPNhT/I8
T07M6lUeOywWHRGtK3K+0plJCTRC9WINUvkVeT9iUWZFQJaLBCg8Sy7EhBcDcv3z
REESVfstGuaQSVdhHhyq+fwQObt4OTp8v5vhqfyg7nRS+uzW7ZlWTiPSO1OPy5ZD
xjW7Yymq0aAjXeBUUjgdnWd+oSDR7PElvPoWJWm6/Lra8NGhrMDRS02Camh913r1
1BPEQGVBaWfokCTmIlHXBDpxqwl1Kw/BSXmHfNph0iWnilZE1AoH3LcnyWsx3ca8
sodQYCXXMbZ0RteckLW0o0rSK6oFZTOWTFT6gO2cFEytKwZgZcYhw/8caLFxw+ND
5e5e2jeZGejGm+sjhqQpbyIMxuP/8QNAsvuP/eE6HE1isTsOmIi32GIYN2u5J1ii
BexLZ67yYMteW0N6JovywZC93wVf9qYANNaQg/4fYLOc1zgLgFNDXeXGsv4V0F6b
ENkVRLXAo1lfFPiAPx49h0p9HDmFLBaSuW7tZC1o7g1G38wC26Mp9d1bRBBpaGoc
Ec02rCtr6VzdzS/0KqCgJylg11doSpMfDsasFIWzxmBpHnM7OXqirxOeV1wUwydL
fuI+/ba7lP/EY80rHFw5cimFGwgD9qzMHAyJOj7vM13vmHSa3wP7wtYEQbWQlACQ
2OCKbQuTAXXN1tuLEmDClJiNc8FIozGmUmHYS4X3E5kXThLk398dVWn5W/9Jr6Ut
pHGPMCAqoa3znUkvD5jthcxfJTlGY2HOrQqbq5u7a9hZCyL/w2RxulzcTLGI0H3h
28qnT/Y1xzqTQgr5U4+TXcXTjuJPkhfZEw9FkBJOYy34X2TEHPk1Ag1C0gdtWXco
J8CGDAre1F79ZDv2td8uzLPsJ8TU2T3LRzGpRATXf+z7c4nTo6BjYzPwNKfBhb9l
6OoQnl03R9N41aG+SR8aBdYWoi62r1xKvabKHQHfN3pHWkPPuKRyzYroEZSC4/Xc
2RbfgVKpKo+EpOVNgk/BT0vnPxoxgD2fv2ORHQPR12LFzqUT4EPKZ/5ObScHhO+F
y7soQEFLPo35mdqUeTM1BV1O1tTbjDDvLV86P/vtXKmwuRHHKF5pYm2CNBtUi6s2
Dvzrn01ACRJHCgnTRnprbN9i8bfVS2DV5mX2tabcb0FDEymcVYpLq8xVdYhbI0rb
6iw29JmDEMncyLEfswBrWZCAVmtZCH08FzCU1z0UsVCF5Y8IHWDEYwXt9XJwCrCy
TcLlxS1n0xfYaiATXLIArOL0r6FVmmRhnziV9fyXd/m/yxAkOAWMe4YdrALz40D3
hBL0eE084XtR2Nn4H1K9nE5yzSYGReI7gsr54K782cBNeV0CXDosvqx+pAC6hIQ1
IhqZMqZfzMQvDe5uuuy75hfBLfi/X9vQg/ntiC7wOdjFACnT7UtE2cUSj/QTil9u
jFsZsZJynmMbozhvCUmhgzoMqzcxaLykFScmH9/ZmIJ3R3iUId9m+3m52H9lgkvU
HnwFkLiEkfApkQ2736bLHPf3UAn7MgWQk2NMsobTU2E=
`pragma protect end_protected
