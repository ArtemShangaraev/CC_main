// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:32:40 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
by4y+ssvIok223cdnBQu/3PXiyJkd+eZwH+bPUgzd5BKKNfnQeIrAg4f7YtCdge1
dhsoD0/e5itR2tO5sZBjzKAQ7cy1otAwAmAXkUkU7HEGztZcopUD84dgNG0x/1GT
gnPpSHuSxMuHkPqWiUuTaWeGBPpHeJgV1MJffCmQi+c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
X/geykMR7mzSqSz97lAXair3TiqZ4fs7ZDW0QJmWcPxGonRKvJEDyFlWcUPk0PQ9
uFxopsbfzBnfbUvWnpnFZKTRop9MmPDisXk1+MXtJEV3QBaR7xPEy2d/f3o9vZdG
g4ILbhPIg6OQU3tW19jJ/fl83fdUn64os41WEkWgNRE3GKjZBjVKZY3vNA/la3Tb
ZAMGXuM9hG9AAVkgkgLKNjA5YzvN3pTjCw/soCOc0UfpVtKbABf9JiS6Ke2jDLk/
hF1FDgcCcBzMklgU50NymG0kGIyrZ3ZoOd+e0XE/fHpIzWSTQDlRdJ6uC4cnE6T7
vNZ2GDMEJ4MvdAAlrwCwrP/dMx0cUJWCX1XFOyc/Wxtk9+HV80r4RZG23dbttCyw
8Mg0MrqO2IbW+I+LxyjArLh8xg5g8wx54/jp1BKAPvlsVwO9vbuUhGSV5Dn31cvS
265LY04HJNhXSGP3vkAuj4Yk29DFLaH1WYCVHTbY/H4W72qf4xZi0oSvjQ6hjA3m
WyHX135rrrYwEaOA9WqhaUhagSIEhQbNQk2MgXFNZOYuKtsHb0pbkDLayuZDon65
5IplDyON6PMM+L//zXoCcU6Bq07E5ao3Ww4RaxQkiKOSKvAE7eHfkIatGpukFHpa
+/4yHIhbPXmTG/LgMUL3P3dcKob3q02BkogunLzxoGdXi77rsoMq7JQbxE1J0A6o
+vAomSNvmAV3blqKoONwj75HMVbb80mhjv0gPcGfjawS1JsFmzoAXRpLFBCaCORE
UvPisIsvxrCwSeWw1wbuwgsNgPSiDHinTwxC12CnjgJojh8pEDEfMIyIsjlIN8GA
/aO5AF2WHn1fODQXsZOUcRZfsudJIZ1CIzoiUCPLjh4Ft776YFwV3Kw1rNMDGs9h
gjDicXuoaaRUVEcDUJB/q+HRYhuIhcKiZxIWf21zwpvJl6bd+VN1VQ4IGbjvjdKR
e7lhVytksSxPWq3QOliXfBkolrJ0PD+GObn+GBonygNek/XgAEzCqPiQ0+hE+gYl
WtMv7vCzaGKdB2kbI+AYMU4CG1UdM6H6AdLXp1PXAupvqZrFQBdLf2kXbaT4tYCk
Qfv+olCjpT+w7kXimLbx4c5ysPGZ87Uii39CDG8b6bGL1J4YOPVOXSJu/oP2l20k
AbfJh6xdl+Ol5+dqxH4/DkCBxGnjXc+QtEyRd1VnOq0sLqRiLkzRk8cD8+Uw0eQM
uz1ATthwsTC5mhuDh5MoViiPhZkp2inB/0Q4RXMjaK+gY6e959UyqOyFActah563
8KW7wjzRGCy04K+NxZIsbZnZhtb7F5BCZ4+8ZodJV31YtXLsrKy8VwLzhvQch6As
WlAPoptoRX4iH8MS0p3SERnw8Wi7Z2s1Ga2dTkA3353Qgk0NkBoRZV9w4JQ689cT
bZi1eC68xSp3yQdgYkgjTSgBCqDRXsGOVABKtuP82ZdpFWSGhPCXRLDP5AtM/zQp
dYUCq1W/q8Ipm9wJT09i8hjATNoBKfSj/YBBbccJwAsNnpRSoNhmPAH/nXcwv1gq
DlgUKzJqpFrolNQRU+ppC4+QZqS2hyVECaP5kso3Ye/c9Uglok9Tg5Z6qfVup3Gm
Qrh3NUO5laOU1kXRtQYuwg88CK02TQjW8T0IwfwZTPg9gzOZiLR8R1c5HrBFidbd
+25t+mdCihx610PLlE1P0MVKvgMmaFqxHm6qdnPOUG/JdIzOEg78Bgr15B+i8by1
rnpGmgwT6PTfSb17Gys2vaGP8CL2OUNjn/DTjpxiQrC+ssgrkP04GNzqSOhmrsIn
Q4i45ulIscMRQyo0rG5x0gXqLne4TG4nw4EzcxY/ONS38pV4/gWAMlS9tK/pR44j
nwiMvLpXo1NgN6or4UUT8y8sjL7F9dFh+8Taaij6BRnkh3BpJnwauYHuHvptanc9
aQyYCl7tSySEP2kiT2BixmGiM3m6IuHzdy8Ss7FvOURdAgQKQVMOHOYZAoaaRNK1
SpI5OKQ9miOAaAhHdVYZ6Fh4TUqyHNE6nGj31VFPXWC3BTK4allmef4ifrrh/26+
imZA3OtVuUz27K+LqEnYAU8/o3LFLGmFDZt6AfASr2r6AFO60350ZzfiqgWThwJP
qxFTb/+v4EkFDSjU/5INVjwihZm3fiMlRtSEvMe+IaOQCy2J9mwTTK9qA3xvvDRZ
ZpmaDc6kphkMxA6hKHCOZ7KmCF2w6wSimwP99l0Yg693f+bpL+fLXvVMYjZQBpRJ
D/ZbwmbWMPmYQEdfUv4AZBoGkx5gMcuM2vycCGK2w1vL9I0H9pOeWIBbfSMmVzJc
oSStPEzwx2IFaOpolCGr7ll+9dcMJMkIQumgx2eWlxGRn0agZRAd2ZMrvWlx6bBn
DIauBXf8XFbInszO3hOmfUL+W4ItkGYP5z9KmMsE78R9ktf3Sd/NafO2Z70s6R+N
BOYgb01GVeQaYLXNscP9stl3Ig1cSKd5AZw6Bk0FZh5A2qMJIcWItXMNuTeG13ho
rDg2Ou+PBlh1MLZw6RNaLZ+J6DEUjHAqNpJIAEsyRHdeVSU7rw+SMvwbe7ZFk+ts
T55jhbAHi3CNitZ7LgaYzyRxZRopwufw4zys/UkyofhiMuc/o610dM4bIIRgieKI
706YoVliX3KmkgbmNC495yagDPLA9VyEPY2rRllvPJPhH6o3dwN6o8f5K0p/h2J3
KFD74Wp+OS4iLq85IFY1OUEgY9MnuNiSqKsg/POcjnfYROdins9ODhwnWqGj1s2Q
ZgYc+9qKyB2i3JJRpqFthk4MPWOLwH9UmmdOPs9lHu0psVDH0AzhpDGm6WsqGh8V
R3vjHRK6x8h+dCeq1WMeGxD+EXzbe5prd/e0DnSfdX6q0CvPU197puRF/h2+CzJ0
YqhEr9wzs4M7uGamoSXK0XA1al1FBFtTNqXz2MnCH27b8qwtk+SyiL45B+76SsDh
b9kyr5/6KxZF683Z9zRtJKHPHgUGU/QLvGx2TBAm/S1QhzXsfDkEoNQ1OcShuchO
tQeqM0fjiGwFeieMF68tQfbcZVRmbgSdDEDj8gHtz3wUm+AO7y3j3ScrvfRF4XP7
ahVyYoQZUnF8wC4RXHFvWDU//jaTHBhWsnSwaW8OHIz16rtazTXBA0axx+Xx2nQM
sOiXsFEgEHV9fG8Al9JG+h8ad8kNdUz3R5hHNS5wQZFFgTfl7kdS/BFzTcUot+Gp
jV6+NkEA2CPhtO2tIgIB5XuwWSh36+UalwQ3uXy2Ucarorv3TQiRC4auvujm1auK
PY7+cYi2V1o1PVzBA2kbsjmbpsgesir+aickOUjoh1hvS6IgfLl0gdDvoRcyMMWI
n7/coWN8rOy3OArXtyjABrIHvc8aoVWEcd1eKMZDsUNwnikA6rvPt+0ct/ms46kV
X2AgihVv4UTiP5FAxd/Q2FBVuaJ1aLkRkUNn8KBAIW85SvF/QxHkch3notg3joua
uYFuyOr8QrzDpBL1o/nSA+EZ3DAEGnyeZZRDIOROgJx6sjQXvZHUQbbHYTdhXNLr
a3dOE/dZHtv5d6u+UzLqj0gtWL0ThrrYKpo2ocGzcVU0ORENEZMolHEAP6ywmHtY
uPlkTYTJ+sMoZzAKal+ygnMUPa+3nN1RzTxx38ilGqueBIEcoDEioPj/gFRavOQT
chEEzki8/pyvu78o3+/qFefz5i6FwC4nBy3pJ75M1j2IHeelB8AlstxyHCqm6y56
zXkfk3j3Kc63jjlxAHwTBRtsqguL2/aXRxzEvOKJ4mXPxC1SrnGHNHDwhq+cpeZC
u8o655/TehYlTTCT/bd7/ygRX6KXBtU3BWtbB7RZ5rjLT7JDnoy7l/y1USNAvihZ
7QRyl3zALeqHQs3vSkbJjigjhtY5psbHzhxwZ/NM+VU3TQ3H1vUjRxSFq+YuTteK
MQ/qlTSMVzTehH3L/m/iGTtaLm6hbpsPuvsjQY2sbngvtvj7IQpHgcS7UGSAtTKC
FJ628KM0Yi73ZoMu9jRLnjrt5FtUvYkQEMC3vVGCFucx2NO9YIMH1fN/YHWYsuVp
ZZdHlWYwSAmqFdu054/1NBysLVY4Z8N37ndr7djyR/T/6MrJv/AUuXdsll6zxuY1
ymrchDLTPFatxBPkQFzUNp/zUP31344tQ7xapXq/85OZdxaYGrLCxOA8WDtvm1xe
Bq7seUDKmhADd/ktCqzzlKKjmJt1s9folUIDVJlRe6YFQU1stN6Av/t9OQdl6pnd
IkoN6d3RwZ2sfWQFqX8i3mNaz6nLnC0yM+GprWlb29AA8a+5IwRcd6Zbc/2CKYs/
T/RIh59hUYmzZ6+iH5VZaHoteFt7IXwJaymJDCf7KVNnGaQVoLCPajQ+Hnml3ybq
A+pGE4fcrEI7cvkPqzffOaincT/yUHY7EfM1oRyCbUDi+KurzMmyzQvskoA9SAVD
qdOZyRwectqLx4XAPqIKjyM50r7w8WxBKpQBBYLRAMdSzzH0vdFDWgzRj5WzMMaD
+v0jcUXCh9oiRRil6BJnZGeMNLwGudNPqKZ+6Ut3oItWWOHO5q/MNzhWPPe9XWHD
v3ouGWaMkdQC4LOjwmCFvkwjxx6imh7uSGeS2ETEJTvawuU5f6Lib9qpZUJFg7ts
NcnoupYiQQvYdl/Zs2iEe0t+yYsw9FGPvMWJyPC6i2f/RZJtPwRiWjCtxQ4BCh0T
z0qe0bDYGzrGWO4jtiRni4EsLDOXF6UgrYR2GdfchPq5TGB2lYQLYqkjeRll8nZ8
g/2U9n22muexWIHhmH27s/uwJ10H2jpVxIW2l/PrbTfS+NzSThuTV6LOueAmn4Tr
bF+2ePqKAuuulMPGPUavvhjZYVqHnIxTeORnYFJwRiOJ8gTv+3lrfIFof9Y+PGED
/I9HUMygDrmbLY7VPgBdc0ODMzkT40q7yCmKySB2TVVZCwWUIAi57nn5aDk7WHus
xld4RYFfRCgs6IaKWdC84nAL381jgZ2Qezbv4qU7Ztm7rmsO+4YlEedfl32DDKqj
kQBx1ZoLp2AcM5+Wp8mb63ToHm7u+6Czv8VoYtSaIQbJjgjuoL7ZKyhGyC+HxirJ
rQa9TR3aCz14SDk7zk3sS8+j4vn+CiYO3UweK1jFT9bIHFyFmUC263UjxL0vDLOV
9cvjZZwMK/UW1EjjRERz6c3ptreGivrbYwpjfa43HagZy5FbNzntTkvlXu+JIWXK
d6Dp3ObIDlIbleqHXOzPdLSv2LWmfAkCt8PNtcEIM0k5ixU/6SDMcRQKj3S0kumR
BlgJ/NGG6dykIw0/7rnqbQqDXyOImC99UjC26nhsrFNgefDsWsqv7YNeq2cU1xL7
jT4sfe9VcVWVad0b7DZ1aUoZb0lDuS7gsPLHJYwlIBlowMAUrSgIuzOIl+ICZuW3
KZS68wDGMtiDPlmeGZDlx6fIdIjlAjdNF1M1eHoOsVslRU/QHKfUskZrbOJ/TYwR
PXexDgG/AiddU1k+mttYBXwnNwvWEemZfJmug/WQedMEZ+3oYgbgYL9ZEAgdWmaG
So8mz/Z7W0439a3yAatcDsHFs4pp6WvADweHhztUf1t1ZCUansfgunGbmChQA2M0
iWjPv7iU0vuc4EGBNl6WYYQfPxp4JmDf3GdZmlVPMdppJxwxejpNyJ1hfdPPr8hO
25WOxvN2hjPrI5frKaeEgoRepNejPZNpcoM5EIW3rbPqHZXJjZnwq4Ao5AE7dNd7
iKfl+zCooT8e5L0r29/IzKVLkm5Pz9LktolqNEkC4PH5fQV++SjTCml6acfa2QMH
kQsRBi2jb+NTzEe0FM9te+2YmzJDuBu0zqxbJqD8f8oZvImWRjCJPH1wvXBmcMfP
hfc+wUj+OsJlMUv2Wz9/iAix0N1n099kzDTOQxJC8mUAc/OWdMsqx8mFBxopwgr4
EZ2qKQh/WfR2Y1dRLhCajsAcMMQxvrHzZ4UzCw9hVyXZyrFBHIq/iwvoXQGO4ekT
fQ7Ng4CkiBPvk4MLw5ASdlVbhkzVcsDZUEwZmqzXq+x3IulOc5QcnTcqWxUdFq8z
OYnzDCRMbhk0MYvw74eo1xkKPDmgUJ1eQzlvcm51139b4GhFIt+6XMR7ELzkorWS
usR0SbKvJoeofADdcDioyibKviyUlHOTCPgHVfbBeQk5vZfC7/OWN5KEW3XsTrWB
vv19jiWoqQx68KGIIhdc3xpLLFEx4RaigaXsu453SiLcMdOJ5tyRrTafhnYE1I9N
Law+GKn22aipJt6SjPNZICVfmRj8NNp3hhyHt4sQgXNLjKL7CiNgeGjZVESEm26G
fza0IMFCGktLk/WkNaFL7u7x21/YFhSWp9padwiAQaUscN5IrdMePKjKMBTrLfOw
63OfATRfvldxJW4Ju2ssonSCL/f6IF6cc7V58itSKTPraEHXqG/Ens6VBUTHc+2p
/vhkfyCakgv4BkuhXGsYypatWCPLUbS74+ABTDOY9XmQIDOUuh7KsoAfORhfJhgg
DUh+fTaXK7DXrczzAY5jF8AguhOGOed+iA7A3LxEoUhobCdPRbAtCAgRGNTTSktV
iL/cr3nT61iTc/lig5sP52Sii9stNTpJ0rW2+fkdg2qGuwaiPlgupcOVwALnNIpE
5+LhhaK98Rcd5WYRaX6YwDo6kiRvaPsCngLBXTP5RM0ZTDkydOKczzwH/6d2ItFN
YcuozOdm+uYzYDYExI1HwuTZGv1ITup6UudjRgyeAdoUTYfxenZnJs1qcQxlPYA5
86zSbCR29xbSO/iwJALYRpd/qayeGUzuy/SiE/Rj42GaBBIZCv51E6EQYeuyb9YY
cuEGETYi1YKhIiN14sq6LeNqtz3T8xPrkmIeNe2Vp6NZfDd4/J2d7a4TzuAtbLhT
oHuOiYmZO5hNLz2NzndAcLv/j4xvdBRkjpYTE8/NHvn4sr7o/Z2XlXSf1MW9Owxq
IneGX8uwnkgi9pvsPNGiC9egrtzhnHO9wJnHMeMUWLMuv0fbYipl554ooAV8iAEQ
mACVpU+Smk5NOid6Vb/43goZbBZBoL2v2S6A5TY3ZeKWy6SSr/DxYsIMLfKjr+J1
LRPkTvX+hnREdvrxlBbhd2fePdrBLstLkecr6CpCz4+wRV9I/czdZU+YOp1bZxuD
VlY7qp1yAKxv9av10NS3zkSvQaBoXdXcpzaC1SoM9ndICDFQGu1ZNabuFKX/bGF4
c4RSDfoSshjA8XTHa57bBkiFkzdOcqGjzXGEI7h5xbrGBw/6CFBZk7fYttXnsSbq
qV9QXgDDGGIQ6L9c05iWkjP0+PiqG+suixNgG/GxSh1Ve2C4X4SHaap0FU5quZHX
M0xQAyhy9JntMHka23xikaP7XuGSRZXQz/AyapeQXA+uI5EASJWdicZvDMBcRcaI
FGHBuDgxwEOxv3TkF4ekj9CoUFLgrRqLygxrBvnGDWEDU06WNjAWmFqmCeTtvSOj
0YC1cBVFwvb3teMlWQ44Q/dgjzQdsF4Q/WFYPta1OTDblqYxohgLmE4d3STcVFZy
0b+WvL4o2BH6bov6MdCkl13HgA5/Q9ZibEoHw97mzxxAr2+3F1Ex8AIHyr4Qg5xS
DppLy5fbtIVHYI1BuT9IO8DpYHmIbMMpoPlO4T2onQrOzsq1uLK9h1MXquuhx8Xz
xun0i7W5ytCcmyfFAfllDs8pxDcnloZqORKRomqgi+k5B9CGglcoEFSDYLhyOVRn
7GIMaqipWl0tYPDVPB/EKArdN11GoPrrJFkq10P7A8f975iWBOfftCJO04Akfiem
3iO9Zthj7OLIbalUAjOhaun40ofyrfaoEdbjeP2ux/X47Y0Q9iLFCDItTU5CowrE
XYg5m/xH1zQWECdflI1EBWICT8+EsH3ACq7z+pgh9eRewmTfQDe+cqmeHhJ1Hg5g
U3sCNLuk2jKZmWzT1n3PNMliBUdx4o4G+TEmsuociUmMqc5pjC09XYrOR1wE4h2F
BjhChRTjv4C9XgFu8WLxKpiKAoJZZCU1ryKj7CMioSQdrURaGSFRnKbIwexYzf0u
Sh36HXvJDfpgmDLiQq2CRU9LzF6DmNevGdGTnXC9YOLp7Z/GbEY9U2fpQBqnKh0k
blVRDv7qLz0xKo1Ia28507mt2OQvBQxQ3vvpehZiBQ8c2Q+xAx7Jssj/bmuieq1W
hVvVl6OAxUvObBfzLAPs9QGxjSRzHWtoci8YjuwdGoX64OxiQEVOB1sf0KqKf5Bg
Y0Rs7x+qol8OYg19StfRdabmsvNdFkPHJ/7HeKWUBD5n6T87QsAwuIDpLiuPC1tm
Ql2n1VmQBgKLr9bN22dW1JezTsyW8VNviGd3ZCqSBKdYxlW7p1nlyvFAnpw18aD4
byiem7WSW65RQHm3N/KOasv+X26LkNelJ2SHIG8nT2l59NwYKpVc/95vzOVVZ0CX
eSkf7YgZFjJVcufbCUco9OXZVrJrF6pUzQZfJlj0cD27CPkqjP3sdqwFbvMLgjbF
Poq63emxKAaYJjSsMVT4m+FzDMa1w1253IWQjx+zcz0DHhD89oQe6cbTNL+eOjat
qWgEhmxuogqOg26co/cT9UlHUjMcfwSi96H4BMPX6EQ/zeAq6ifM8Ep7cQCKBbAR
b6wEJtTbKQ1ONgvGw0oEOzkvnok3Vs0j4m63KGAkw0HBj8u1Wd2tXD2233YoaUhi
HteTdML0uJG9QktDBRbOrJWzWztqAUOPIUl6tBVWXvd2FF8Y6o993HYYp+U5KpWg
ZMROjJz72WqijJIYSCTg/ygpHSAuhYPCVMMaVd2CjrihS9gxI2TdTuKcrVYvS7ce
IG53aEiN9W+dwKsAZYNO3WqkJ4w4CLcpvQ+rlY3DA8ktj02w7T6+P9g63zt2bRlg
yIlmkMicQ8PsHcSduRgqn8k7IIYhT6VBJ/dYjVYWOVrpat9ar6rVHPewJBLDnBeM
hOp+zB1TsmnvKR72zz9uMICNsCe7qLrh48ZPp+4mMCvoo6RyXm2LlY8X/XjVNh7Y
BUyAos4DOoxQQS8CqC467xvcEc5tc2+MmfJvFuFZO60taQsZaskGtak4JEQUHJMi
aCWaL/GMknvCgEpLF9Hr08ygz0bcDy120zRjZh1+qhrg3ymgq6FmNB07T1gVmlfu
vfHly028p95SVVb9vfOF1gYBPnMR0wMju9ZEATluORnDzaMegLkbDvLLq8CM3KVz
yekwJaWbDCD7w+mr+y7NfLCrlDEXTJqIzXRz5UbHy3WJNr7DMKyGcrklR9qFMMtp
xq2VeDB0g77qQQl/cXO2ZZmnBX4jE5/QRJ7KWyb3uN4OabT5Vro25xTMx0HR8Lkr
YXU5bJYvhqSlQe49yUYml8pGmL6oilr0f5uViGrDrFNOtxDMvtDQgFrP5DPvlTMb
AcKVDngxMK2bJdbV3S5FxWmAUj/YQL5cOGmTne2SqC/Y+EU4Oro6G31NfuaY413N
7oxaN/1LRf9noSRIEizFkP/nnHV6HA2p17TPt8sLl0MF10jqofXbc4tV5d/LLuC9
aRBhxa9Zef33dnqyqHbDOFBMDnP5URm2YP/Tw+Np0hH+X+JyDF8FCiTLNVqSFWSp
1tO+7ajXVx9btBZQUjftQ0UfXdRNwOs7euJY5IUqj/oCZJ4R+o0nS95yCO4TbW+r
54zwGWJoRIuGHbtCpuZJ6cIk42yJ9WCtMd/Po3vY65WIMfrV/lNH572Zaw8YrdJp
0zKz1nHcoZRW4r7D45RYNp/2BYmOX9cmGOJlxBlWe3CR8QwqXopKTAM3v2RkXUXj
qUxblZi281lUEnd2Yf+R7PzOtAK2faNrdBNXXJklr76M+D5zgdokPnggfMdR0nsK
E3yHQe2uepqkMoACNxDvIS39Ur4XIGRJ6PXys1kHr/EJJecNkFVz1Wg5syaX7rWo
UgYWYC5bNoKlHzh2LmykghSsUjTagbUrcScV8EGuEljaaw0CgUehcCLP0B1NFgIG
RRx9RRG8e4hB25We2ppMIzaYpiV1gaqqL5BwyNEXdAflVUSp1hzNbFn2h3EfWab0
YiTmHaaDel+Xdzs11jX/b5hV6UEKixx3BELPdzqrZqvaKIxwWykaBkzN4jh9sTix
Fv50G1Gnm5zxshqA1V/VfI35qREpL+AgVIwir2PnpRAESIgPgusIU4zxzVmDrl3P
ILZCmUu6GMFq2+8iYjay1XW2JWum+86OSOsyABdpn/6OMjGVKQKoOV70V6HnUFfg
Ok1sodZtTMxDxB82Bdi55a99FtcIVojAGxfIl4Gr1kAlNarB6ZtcWWTBG+4/nUfQ
wKtfeVjCOqdgK01oPDuLX2yKaiCbKriPKLra34WVVSQYFMAy9YvX4abo1IvbDNkL
Cp+8tIMsu8Ysu7ap2HmmX26gCWYB/6lHnwPuXjqBH+u6uCQZc/e5IEXUTDw2T19A
NmBc5rCHcOCt/nKy94Sf/IDl5zTGfOVU1Su7MxEgdEE3ZuYX0+YIXLswPTCtCb7w
EWpwooY1BtatD5hjgqoovNiLXT4lsLY+Dro4BAOcbMCRDHQvkx12r831dOYV3J2E
t/uIVr0MARNmfxRqt6ScVbBwg4NtLSmh76roFR4p0NRcu+neTbCK0+19tnnDXcW6
vT5g9oNHShCLutEt2IW+V1c0+qxoUc8VjyYpu2nFXAHnX24zWt2EDrrIye3INcf4
7/fkYanhtWRa5i/svB+rABMDl/klqgLltVkB+lJVWoQ14ukjiV2XWm4JXoWz7ctw
azMHbY4NoRUESLXBAgpLG34xUhcW+aDcIooN56JqWaG2DhMn0vUPYikdfgToceVd
IK7jf4jZCoOUgdI6Ew5xxJWIgtzVeAEHF3qEO3ZhLt4cWgWCFvoLkc3D9eybBenl
X3fsM6c95y6XWsqOHl2NZZ4TiaUWcPuZyklMTzVjBre2igCHJGow00jhei2P3I6/
JPasMQGfuTnh6QfO/iIvYEaukNRYnGL1ksYIAp0YikPijfxcfM/XLcvnbOwe/Jgt
8PdcKnNghA5z+ph0wDzCT4YnWf5nAAbqvVmkGQ2vzS6AQ/T8ry9SdwRVkDyZtmQT
nB/41+TiGQOQ4q1jaJ2mEWQq0Py/J4t0eSQaCRifUeRpXR2p6mfOsbHHDiGsuiDw
I+Ccl7uYI6thi8QsAgRutbFjfBPvDZL4enMyuYoF2cxYmB7n1bE2oZMD6AAIizqM
iwqGt/ZhCjW0snmy03naBGKE7FWjiCnoLpxrqqfbw63CgEYzSfSUY0Qyo5Eco+4w
6fWukBCBk74UyjYdwZL15s/2WocegrnQnQIfe5kWTByNaurAnQvl3DljdhruP8fM
5FrqxfFn/bnDnFIgwrMmeji98O3Ek7hB27/3HTNFrHjHGZh/qiowh/HIrB/C2gxp
vQmeV7yhxORCRv3YlqAAbOA5/UHGNNgpfzdtVTIMKX/0cH4G37wug9f6Cvsn0GEM
FPyCGUywzS6D8MeXWbt4gLdMKG07HWoI1Fhm3gIlNl611Dx6SZj0vE1pBPBv3vr+
w8r4DiEMxZ8Y/bBW+/7X3JdNjy9eDGAVr0CiZQejy5ZhDEGglTcS+/2IuzhnKMMz
Ap90Jhl9nWwhpCk+BWE+iU078AqrS0JFdtz6IVN2Lw3W+O9sFhR0h2kAOEfb32JU
Mf/cI6pjxqpkpkoBXhBnIcf0VnL0TuQMTD2VdJhEnS3XDjCHUNnsqrmdqQFbh+MT
GC9oCr0rYR9jnI1Y7P+Tf4bs+gEDv4+P1VDAtMFvLvqBOBCXmoaCq51xpWEoQRBr
fG0weSiqd7SN6icQHMgslcxvkEnkAFzS5u2LVlfhvX3F/OC8N90mik44Oh1qkWv8
gt2kVYKz51MI4TPRlzYKmNvbympZk+PVCU+LR+tfZKFRomH/NBGjRjUu09QGQjk8
50q7TwrT2gqn7RNX04o2TeOUvsKE8Ff+0/IjB+P0kY34BXUXr4HQtIV3HDQjM+aU
io2omnUJjxW00MiLYNKZb1ClRl8TkfRnycAbOYTBT4RLT3j6/GWuIdhfApuHgu8Q
rg364Lt0YQ8rVbrJf4muVUik2u30bZJyXqm3KfGcwlcJVpIPLTcM9kuytgXipkWu
A0ohguizLSsfhMmD62NbQYXZ2YLamaKfx3yG9Euo8ZlIPutRFqRJ5+/ep+f+vN6W
Jm+tsq1lxttV8h6REYzN4gmR6Qz7+DpJiGX5/M44OpqpEOjVT0+wLiHMGIqhxTgc
rLw0aSbApWBdS7nuLySUOxHkS0cv8MNe3X+nniAH2hL/D05ow7xzCPXxAVQtRRpE
KCRZ2+q4Ra9RPaHAAP2L0VCu0COBQu08ATs9IGRtOXhghX7M4pDEJ2oiIT1TmgfG
T2wdTLynk6QuUUsQVZLYNzG9bIOr63bYTeuCHJgExjEOK1Og69xFd7Q7WfgsccRQ
cS0vSsd6Ssflwy8UUi2ckGGw6C/r/HYWFC59+DanA84AEqbG5+mUW0abPvev7yR1
y/IymawY/9yDxsoU3b3fRouu7ooUSwOOykUEl6g3Zx7cPCOPB5vO/Be2ojp4Jo7O
uKfd6Xrg18IQnmaaDuWVecZvI5NiEuungDe3cCqUIH9NAZgG6s4Wmm5ddK8pvRLA
ain7RT4gIDWZUNTEuNisip0REmV6G9VlUgEqAHJeXy7apaFJztTTrWxMFzIDtWsb
llSCLi02RtOo8KsNaoelNbEMKxkEy/7v9PXGftubiD1OYxHqI8tge6DW403q/XnX
VUKhnIcnskJCsQbSzgo78ZoYL0IkgXOOzpogIgrjyzWumXapfDQnM8KUSXj86SSG
NiV4NfoCbUdYdsM/Y5C5+LRhSeW8mCpRHZKjb75mI3b5++TNPmtrynKANLjPNk6z
5DIRRXnS2xP4cfynxKHfO3cfxrd+rv8fJz2Wel0oxFMVNo8y2iiVciFqgnkUGJtO
9i45TgdVv1sUzU4VeQJIeKFBIrwaiwROfXAWw75aelRzI9R30USvPzp4fE9gOXQn
LrhUsZPinTYF8PAOtT+Lfk9xZVYJgUNa70n3vpeM/FEhQoSUen5ILbmuPONArWCu
pmK2JgSDCCb8+K6K5Wbc4u6pWoDYfHBUy3jXIHnvF9/ZQSYjcfI8sVwNrMXjfM2y
KYuHcPMXjSkGRpLCuHfz385dH8AARtOhYzPaTkmrnzColpnTGI0uJOxSHzG3J07i
`pragma protect end_protected
